`timescale 1 ns/100 ps
// Version: v11.6 11.6.0.34


module COREAHBLITE_SLAVEARBITER_slave_arbiter_4(
       masterAddrInProg_i_2,
       N_290,
       N_63,
       CoreAHBLite_0_AHBmslave5_HREADY_i_0,
       un1_masterAddrInProg_6,
       N_387,
       N_259,
       N_368,
       N_408,
       N_283,
       N_409,
       N_284,
       N_5,
       N_282,
       N_342,
       N_293,
       N_341,
       N_292,
       N_340,
       N_291,
       FAB_CLK,
       crc_ahb_ip_MSS_0_M2F_RESET_N
    );
output [0:0] masterAddrInProg_i_2;
input  N_290;
input  N_63;
input  CoreAHBLite_0_AHBmslave5_HREADY_i_0;
output un1_masterAddrInProg_6;
output N_387;
input  N_259;
input  N_368;
output N_408;
input  N_283;
output N_409;
input  N_284;
output N_5;
input  N_282;
output N_342;
input  N_293;
output N_341;
input  N_292;
output N_340;
input  N_291;
input  FAB_CLK;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;

    wire \arbRegSMCurrentState_ns_0[1] , 
        \arbRegSMCurrentState[2]_net_1 , N_164, 
        un1_masterAddrInProg_6_0_a2_0_a2_1, \masterAddrInProg_i_0[1] , 
        \masterAddrInProg_i_0[3] , \masterAddrInProg_i_0[2] , 
        \MASTERADDRINPROG_iv_i_0[0] , 
        \MASTERADDRINPROG_iv_i_a4_1_0[0] , 
        \MASTERADDRINPROG_iv_i_a4_0_0[0] , 
        \arbRegSMCurrentState_ns_a4_0_0[2] , 
        \arbRegSMCurrentState[1]_net_1 , N_154, N_187, 
        \arbRegSMCurrentState_ns[2] , N_170, N_169, N_168, 
        \arbRegSMCurrentState[9]_net_1 , 
        \arbRegSMCurrentState[13]_net_1 , 
        \arbRegSMCurrentState[5]_net_1 , \arbRegSMCurrentState_ns[1] , 
        N_163, \arbRegSMCurrentState_ns_2[1] , N_184, N_157, 
        \arbRegSMCurrentState_ns_a4_3_0[1] , 
        \arbRegSMCurrentState[0]_net_1 , N_156, 
        \arbRegSMCurrentState[3]_net_1 , 
        \arbRegSMCurrentState_RNO[0]_net_1 , N_158, 
        \arbRegSMCurrentState_RNO[3]_net_1 , N_160, 
        \arbRegSMCurrentState_RNO[6]_net_1 , 
        \arbRegSMCurrentState_RNO[7]_net_1 , 
        \arbRegSMCurrentState_RNO[10]_net_1 , 
        \arbRegSMCurrentState_RNO[11]_net_1 , 
        \arbRegSMCurrentState_RNO[14]_net_1 , 
        \arbRegSMCurrentState_RNO[15]_net_1 , 
        \arbRegSMCurrentState_ns[13] , 
        \arbRegSMCurrentState[14]_net_1 , \arbRegSMCurrentState_ns[9] , 
        \arbRegSMCurrentState[10]_net_1 , \arbRegSMCurrentState_ns[5] , 
        \arbRegSMCurrentState[6]_net_1 , GND, VCC;
    
    OR3 \arbRegSMCurrentState_RNO[1]  (.A(N_163), .B(
        \arbRegSMCurrentState_ns_0[1] ), .C(
        \arbRegSMCurrentState_ns_2[1] ), .Y(
        \arbRegSMCurrentState_ns[1] ));
    NOR3B \arbRegSMCurrentState_RNIRP91E[0]  (.A(N_259), .B(
        masterAddrInProg_i_2[0]), .C(N_368), .Y(N_387));
    NOR2A \arbRegSMCurrentState_RNI72O91[2]  (.A(N_187), .B(
        \arbRegSMCurrentState[2]_net_1 ), .Y(
        \MASTERADDRINPROG_iv_i_a4_0_0[0] ));
    AO1A \arbRegSMCurrentState_RNO_1[1]  (.A(N_290), .B(
        \arbRegSMCurrentState[2]_net_1 ), .C(N_164), .Y(
        \arbRegSMCurrentState_ns_0[1] ));
    NOR2B \arbRegSMCurrentState_RNI8GFO9[0]  (.A(N_283), .B(
        masterAddrInProg_i_2[0]), .Y(N_408));
    NOR2 \arbRegSMCurrentState_RNIU70V8[0]  (.A(
        \MASTERADDRINPROG_iv_i_0[0] ), .B(N_184), .Y(
        masterAddrInProg_i_2[0]));
    OR2A \arbRegSMCurrentState_RNO[11]  (.A(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .B(
        \masterAddrInProg_i_0[2] ), .Y(
        \arbRegSMCurrentState_RNO[11]_net_1 ));
    DFN1C0 \arbRegSMCurrentState[3]  (.D(
        \arbRegSMCurrentState_RNO[3]_net_1 ), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        \arbRegSMCurrentState[3]_net_1 ));
    OR3 \arbRegSMCurrentState_RNO[2]  (.A(N_170), .B(N_169), .C(N_168), 
        .Y(\arbRegSMCurrentState_ns[2] ));
    OR2A \arbRegSMCurrentState_RNO[7]  (.A(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .B(
        \masterAddrInProg_i_0[1] ), .Y(
        \arbRegSMCurrentState_RNO[7]_net_1 ));
    DFN1C0 \arbRegSMCurrentState[10]  (.D(
        \arbRegSMCurrentState_RNO[10]_net_1 ), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        \arbRegSMCurrentState[10]_net_1 ));
    NOR2A \arbRegSMCurrentState_RNO_0[2]  (.A(
        \arbRegSMCurrentState[3]_net_1 ), .B(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(N_170));
    NOR2A \arbRegSMCurrentState_RNO_4[1]  (.A(
        \arbRegSMCurrentState[1]_net_1 ), .B(N_290), .Y(
        \arbRegSMCurrentState_ns_a4_3_0[1] ));
    NOR3C \arbRegSMCurrentState_RNIH3B41[11]  (.A(
        \masterAddrInProg_i_0[1] ), .B(\masterAddrInProg_i_0[3] ), .C(
        \masterAddrInProg_i_0[2] ), .Y(
        un1_masterAddrInProg_6_0_a2_0_a2_1));
    NOR2A \arbRegSMCurrentState_RNIGNTN9[0]  (.A(
        masterAddrInProg_i_2[0]), .B(N_282), .Y(N_5));
    VCC VCC_i (.Y(VCC));
    NOR3A \arbRegSMCurrentState_RNO_0[1]  (.A(N_154), .B(N_157), .C(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(N_163));
    NOR2B \arbRegSMCurrentState_RNIBSCM9[0]  (.A(N_292), .B(
        masterAddrInProg_i_2[0]), .Y(N_341));
    OA1 \arbRegSMCurrentState_RNO_3[2]  (.A(
        \arbRegSMCurrentState[1]_net_1 ), .B(N_154), .C(N_290), .Y(
        \arbRegSMCurrentState_ns_a4_0_0[2] ));
    NOR2B \arbRegSMCurrentState_RNI9HFO9[0]  (.A(N_284), .B(
        masterAddrInProg_i_2[0]), .Y(N_409));
    OR2B \arbRegSMCurrentState_RNIT6D51[2]  (.A(
        \arbRegSMCurrentState[2]_net_1 ), .B(N_290), .Y(N_156));
    NOR2B \arbRegSMCurrentState_RNO_1[2]  (.A(
        \arbRegSMCurrentState_ns_a4_0_0[2] ), .B(N_63), .Y(N_169));
    OA1A \arbRegSMCurrentState_RNO[0]  (.A(N_158), .B(
        \arbRegSMCurrentState[0]_net_1 ), .C(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(
        \arbRegSMCurrentState_RNO[0]_net_1 ));
    DFN1C0 \arbRegSMCurrentState[0]  (.D(
        \arbRegSMCurrentState_RNO[0]_net_1 ), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        \arbRegSMCurrentState[0]_net_1 ));
    DFN1P0 \arbRegSMCurrentState[7]  (.D(
        \arbRegSMCurrentState_RNO[7]_net_1 ), .CLK(FAB_CLK), .PRE(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(\masterAddrInProg_i_0[1] ));
    OR2A \arbRegSMCurrentState_RNO[15]  (.A(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .B(
        \masterAddrInProg_i_0[3] ), .Y(
        \arbRegSMCurrentState_RNO[15]_net_1 ));
    DFN1C0 \arbRegSMCurrentState[14]  (.D(
        \arbRegSMCurrentState_RNO[14]_net_1 ), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        \arbRegSMCurrentState[14]_net_1 ));
    DFN1C0 \arbRegSMCurrentState[6]  (.D(
        \arbRegSMCurrentState_RNO[6]_net_1 ), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        \arbRegSMCurrentState[6]_net_1 ));
    OA1B \arbRegSMCurrentState_RNO_2[1]  (.A(
        \arbRegSMCurrentState_ns_a4_3_0[1] ), .B(
        \arbRegSMCurrentState[0]_net_1 ), .C(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(
        \arbRegSMCurrentState_ns_2[1] ));
    DFN1C0 \arbRegSMCurrentState[1]  (.D(\arbRegSMCurrentState_ns[1] ), 
        .CLK(FAB_CLK), .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        \arbRegSMCurrentState[1]_net_1 ));
    NOR2 \arbRegSMCurrentState_RNO[6]  (.A(\masterAddrInProg_i_0[1] ), 
        .B(CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(
        \arbRegSMCurrentState_RNO[6]_net_1 ));
    NOR2 \arbRegSMCurrentState_RNO[10]  (.A(\masterAddrInProg_i_0[2] ), 
        .B(CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(
        \arbRegSMCurrentState_RNO[10]_net_1 ));
    NOR3A \arbRegSMCurrentState_RNIASPG2[1]  (.A(N_187), .B(
        \arbRegSMCurrentState[1]_net_1 ), .C(N_154), .Y(
        \MASTERADDRINPROG_iv_i_a4_1_0[0] ));
    AOI1 \arbRegSMCurrentState_RNO_2[2]  (.A(N_63), .B(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .C(N_156), .Y(N_168));
    AO1A \arbRegSMCurrentState_RNO[13]  (.A(N_63), .B(
        \arbRegSMCurrentState[13]_net_1 ), .C(
        \arbRegSMCurrentState[14]_net_1 ), .Y(
        \arbRegSMCurrentState_ns[13] ));
    NOR2A \arbRegSMCurrentState_RNO_3[1]  (.A(
        \arbRegSMCurrentState[1]_net_1 ), .B(N_63), .Y(N_164));
    OR2A \arbRegSMCurrentState_RNO_0[3]  (.A(N_63), .B(N_156), .Y(
        N_160));
    GND GND_i (.Y(GND));
    NOR2 \arbRegSMCurrentState_RNIFMQR[0]  (.A(
        \arbRegSMCurrentState[3]_net_1 ), .B(
        \arbRegSMCurrentState[0]_net_1 ), .Y(N_187));
    MX2 \arbRegSMCurrentState_RNIMP1I4[1]  (.A(
        \MASTERADDRINPROG_iv_i_a4_1_0[0] ), .B(
        \MASTERADDRINPROG_iv_i_a4_0_0[0] ), .S(N_290), .Y(
        \MASTERADDRINPROG_iv_i_0[0] ));
    NOR2B \arbRegSMCurrentState_RNIARCM9[0]  (.A(N_291), .B(
        masterAddrInProg_i_2[0]), .Y(N_340));
    NOR2 \arbRegSMCurrentState_RNO[14]  (.A(\masterAddrInProg_i_0[3] ), 
        .B(CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(
        \arbRegSMCurrentState_RNO[14]_net_1 ));
    DFN1C0 \arbRegSMCurrentState[9]  (.D(\arbRegSMCurrentState_ns[9] ), 
        .CLK(FAB_CLK), .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        \arbRegSMCurrentState[9]_net_1 ));
    DFN1P0 \arbRegSMCurrentState[13]  (.D(
        \arbRegSMCurrentState_ns[13] ), .CLK(FAB_CLK), .PRE(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        \arbRegSMCurrentState[13]_net_1 ));
    DFN1P0 \arbRegSMCurrentState[11]  (.D(
        \arbRegSMCurrentState_RNO[11]_net_1 ), .CLK(FAB_CLK), .PRE(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(\masterAddrInProg_i_0[2] ));
    NOR2A \arbRegSMCurrentState_RNI8EUC4[0]  (.A(N_187), .B(N_63), .Y(
        N_184));
    DFN1C0 \arbRegSMCurrentState[2]  (.D(\arbRegSMCurrentState_ns[2] ), 
        .CLK(FAB_CLK), .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        \arbRegSMCurrentState[2]_net_1 ));
    NOR2A \arbRegSMCurrentState_RNIFBB3A[11]  (.A(
        un1_masterAddrInProg_6_0_a2_0_a2_1), .B(
        masterAddrInProg_i_2[0]), .Y(un1_masterAddrInProg_6));
    OR2A \arbRegSMCurrentState_ns_o2_0[1]  (.A(N_63), .B(N_290), .Y(
        N_157));
    DFN1C0 \arbRegSMCurrentState[5]  (.D(\arbRegSMCurrentState_ns[5] ), 
        .CLK(FAB_CLK), .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        \arbRegSMCurrentState[5]_net_1 ));
    DFN1P0 \arbRegSMCurrentState[15]  (.D(
        \arbRegSMCurrentState_RNO[15]_net_1 ), .CLK(FAB_CLK), .PRE(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(\masterAddrInProg_i_0[3] ));
    AO1D \arbRegSMCurrentState_RNO_0[0]  (.A(N_154), .B(
        \arbRegSMCurrentState[1]_net_1 ), .C(N_157), .Y(N_158));
    AO1A \arbRegSMCurrentState_RNO[5]  (.A(N_63), .B(
        \arbRegSMCurrentState[5]_net_1 ), .C(
        \arbRegSMCurrentState[6]_net_1 ), .Y(
        \arbRegSMCurrentState_ns[5] ));
    NOR2B \arbRegSMCurrentState_RNICTCM9[0]  (.A(N_293), .B(
        masterAddrInProg_i_2[0]), .Y(N_342));
    AO1A \arbRegSMCurrentState_RNO[9]  (.A(N_63), .B(
        \arbRegSMCurrentState[9]_net_1 ), .C(
        \arbRegSMCurrentState[10]_net_1 ), .Y(
        \arbRegSMCurrentState_ns[9] ));
    OA1A \arbRegSMCurrentState_RNO[3]  (.A(N_160), .B(
        \arbRegSMCurrentState[3]_net_1 ), .C(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(
        \arbRegSMCurrentState_RNO[3]_net_1 ));
    OR3 \arbRegSMCurrentState_RNI4R171[13]  (.A(
        \arbRegSMCurrentState[9]_net_1 ), .B(
        \arbRegSMCurrentState[13]_net_1 ), .C(
        \arbRegSMCurrentState[5]_net_1 ), .Y(N_154));
    
endmodule


module COREAHBLITE_SLAVESTAGE_slavestage_5(
       masterDataInProg_0,
       masterAddrInProg_i_2,
       bus_wr_25,
       bus_wr_0,
       bus_wr_1,
       bus_wr_2,
       bus_wr_16,
       bus_wr_3,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA,
       FAB_CLK,
       crc_ahb_ip_MSS_0_M2F_RESET_N,
       CoreAHBLite_0_AHBmslave5_HREADY_i_0,
       N_332,
       N_333,
       N_334,
       N_335,
       N_336,
       N_337,
       N_347,
       N_348,
       N_352,
       N_353,
       N_358,
       N_360,
       N_361,
       N_364,
       N_365,
       N_366,
       N_367,
       N_350,
       N_357,
       N_356,
       N_351,
       N_349,
       N_259,
       regHTRANS,
       masterRegAddrSel,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE,
       regHWRITE,
       defSlaveSMCurrentState_RNIJGOT3,
       m0s5DataSel,
       N_354,
       N_362,
       N_355,
       N_363,
       N_290,
       N_63,
       un1_masterAddrInProg_6,
       N_387,
       N_408,
       N_283,
       N_409,
       N_284,
       N_5,
       N_342,
       N_293,
       N_341,
       N_292,
       N_340,
       N_291
    );
output [0:0] masterDataInProg_0;
output [0:0] masterAddrInProg_i_2;
output bus_wr_25;
output bus_wr_0;
output bus_wr_1;
output bus_wr_2;
output bus_wr_16;
output bus_wr_3;
input  [1:1] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS;
input  [31:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA;
input  FAB_CLK;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;
input  CoreAHBLite_0_AHBmslave5_HREADY_i_0;
output N_332;
output N_333;
output N_334;
output N_335;
output N_336;
output N_337;
output N_347;
output N_348;
output N_352;
output N_353;
output N_358;
output N_360;
output N_361;
output N_364;
output N_365;
output N_366;
output N_367;
output N_350;
output N_357;
output N_356;
output N_351;
output N_349;
output N_259;
input  regHTRANS;
input  masterRegAddrSel;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE;
input  regHWRITE;
input  defSlaveSMCurrentState_RNIJGOT3;
input  m0s5DataSel;
output N_354;
output N_362;
output N_355;
output N_363;
input  N_290;
input  N_63;
output un1_masterAddrInProg_6;
output N_387;
output N_408;
input  N_283;
output N_409;
input  N_284;
output N_5;
output N_342;
input  N_293;
output N_341;
input  N_292;
output N_340;
input  N_291;

    wire \masterDataInProg[0]_net_1 , N_282, N_368, GND, VCC;
    
    NOR2B \masterDataInProg_RNINLG3_13[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[12]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_355));
    DFN1E0C0 \masterDataInProg_0[0]  (.D(masterAddrInProg_i_2[0]), 
        .CLK(FAB_CLK), .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Q(masterDataInProg_0[0])
        );
    NOR2B \masterDataInProg_0_RNI6S7A_3[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[1]), .B(
        masterDataInProg_0[0]), .Y(bus_wr_1));
    NOR2B \masterDataInProg_RNINLG3_6[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[28]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_334));
    NOR2B \masterDataInProg_0_RNI6S7A_2[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[2]), .B(
        masterDataInProg_0[0]), .Y(bus_wr_2));
    NOR2B \masterDataInProg_0_RNI6S7A_8[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[21]), .B(
        masterDataInProg_0[0]), .Y(N_364));
    NOR2B \masterDataInProg_RNINLG3_9[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[23]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_366));
    NOR2B \masterDataInProg_0_RNI6S7A[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[7]), .B(
        masterDataInProg_0[0]), .Y(N_350));
    NOR2B \masterDataInProg_0_RNI6S7A_7[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[22]), .B(
        masterDataInProg_0[0]), .Y(N_365));
    NOR2B \masterDataInProg_0_RNI6S7A_1[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[3]), .B(
        masterDataInProg_0[0]), .Y(bus_wr_3));
    VCC VCC_i (.Y(VCC));
    NOR2B \masterDataInProg_RNINLG3_14[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[11]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_354));
    NOR2B \masterDataInProg_RNINLG3[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[5]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_348));
    NOR2B \masterDataInProg_RNINLG3_0[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[4]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_347));
    NOR2B \masterDataInProg_RNINLG3_2[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[9]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_352));
    NOR2B \masterDataInProg_RNINLG3_4[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[31]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_337));
    NOR2B \masterDataInProg_RNINLG3_5[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[30]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_336));
    NOR2B \masterDataInProg_0_RNI6S7A_6[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[25]), .B(
        masterDataInProg_0[0]), .Y(bus_wr_25));
    NOR2B \masterDataInProg_RNINLG3_1[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[0]), .B(
        \masterDataInProg[0]_net_1 ), .Y(bus_wr_0));
    NOR2B \masterDataInProg_0_RNI6S7A_9[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[20]), .B(
        masterDataInProg_0[0]), .Y(N_363));
    NOR2B \masterDataInProg_0_RNI6S7A_4[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[29]), .B(
        masterDataInProg_0[0]), .Y(N_335));
    DFN1E0C0 \masterDataInProg[0]  (.D(masterAddrInProg_i_2[0]), .CLK(
        FAB_CLK), .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Q(
        \masterDataInProg[0]_net_1 ));
    GND GND_i (.Y(GND));
    NOR2B \masterDataInProg_0_RNI6S7A_14[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[10]), .B(
        masterDataInProg_0[0]), .Y(N_353));
    NOR2B \masterDataInProg_RNINLG3_11[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[16]), .B(
        \masterDataInProg[0]_net_1 ), .Y(bus_wr_16));
    NOR2B \masterDataInProg_RNINLG3_10[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[19]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_362));
    NOR2B \masterDataInProg_0_RNI6S7A_12[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[14]), .B(
        masterDataInProg_0[0]), .Y(N_357));
    NOR2B \masterDataInProg_0_RNI6S7A_0[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[6]), .B(
        masterDataInProg_0[0]), .Y(N_349));
    NOR2 HTRANS_i_0_a2 (.A(defSlaveSMCurrentState_RNIJGOT3), .B(
        m0s5DataSel), .Y(N_368));
    MX2C HWRITE_0_i_0_m2 (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE), .B(regHWRITE), 
        .S(masterRegAddrSel), .Y(N_282));
    NOR2B \masterDataInProg_RNINLG3_8[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[24]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_367));
    COREAHBLITE_SLAVEARBITER_slave_arbiter_4 slave_arbiter (
        .masterAddrInProg_i_2({masterAddrInProg_i_2[0]}), .N_290(N_290)
        , .N_63(N_63), .CoreAHBLite_0_AHBmslave5_HREADY_i_0(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .un1_masterAddrInProg_6(
        un1_masterAddrInProg_6), .N_387(N_387), .N_259(N_259), .N_368(
        N_368), .N_408(N_408), .N_283(N_283), .N_409(N_409), .N_284(
        N_284), .N_5(N_5), .N_282(N_282), .N_342(N_342), .N_293(N_293), 
        .N_341(N_341), .N_292(N_292), .N_340(N_340), .N_291(N_291), 
        .FAB_CLK(FAB_CLK), .crc_ahb_ip_MSS_0_M2F_RESET_N(
        crc_ahb_ip_MSS_0_M2F_RESET_N));
    MX2 HTRANS_i_0_m2 (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS[1]), .B(regHTRANS), 
        .S(masterRegAddrSel), .Y(N_259));
    NOR2B \masterDataInProg_RNINLG3_7[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[27]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_333));
    NOR2B \masterDataInProg_RNINLG3_12[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[15]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_358));
    NOR2B \masterDataInProg_0_RNI6S7A_13[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[13]), .B(
        masterDataInProg_0[0]), .Y(N_356));
    NOR2B \masterDataInProg_0_RNI6S7A_11[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[17]), .B(
        masterDataInProg_0[0]), .Y(N_360));
    NOR2B \masterDataInProg_0_RNI6S7A_10[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[18]), .B(
        masterDataInProg_0[0]), .Y(N_361));
    NOR2B \masterDataInProg_0_RNI6S7A_5[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[26]), .B(
        masterDataInProg_0[0]), .Y(N_332));
    NOR2B \masterDataInProg_RNINLG3_3[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[8]), .B(
        \masterDataInProg[0]_net_1 ), .Y(N_351));
    
endmodule


module COREAHBLITE_DEFAULTSLAVESM_default_slave_sm(
       SDATASELInt,
       N_372,
       N_374,
       defSlaveSMCurrentState_RNI5UNRI,
       N_242,
       defSlaveSMCurrentState_RNIJGOT3,
       N_138,
       N_105_i,
       m0s5DataSel,
       FAB_CLK,
       crc_ahb_ip_MSS_0_M2F_RESET_N
    );
input  [15:6] SDATASELInt;
input  N_372;
input  N_374;
output defSlaveSMCurrentState_RNI5UNRI;
output N_242;
output defSlaveSMCurrentState_RNIJGOT3;
input  N_138;
output N_105_i;
input  m0s5DataSel;
input  FAB_CLK;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;

    wire N_261, N_373, HREADY_M_iv_i_0_i_o2_0, N_339, 
        defSlaveSMNextState_i_a2_0_7_net_1, 
        defSlaveSMNextState_i_a2_0_1_net_1, 
        defSlaveSMNextState_i_a2_0_0_net_1, 
        defSlaveSMNextState_i_a2_0_4_net_1, 
        defSlaveSMNextState_i_a2_0_6_net_1, 
        defSlaveSMNextState_i_a2_0_3_net_1, N_268, 
        defSlaveSMCurrentState_i_0, GND, VCC;
    
    DFN1P0 defSlaveSMCurrentState (.D(defSlaveSMCurrentState_RNIJGOT3), 
        .CLK(FAB_CLK), .PRE(crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(
        defSlaveSMCurrentState_i_0));
    OR2 defSlaveSMCurrentState_RNI5UNRI_inst_1 (.A(N_261), .B(
        HREADY_M_iv_i_0_i_o2_0), .Y(defSlaveSMCurrentState_RNI5UNRI));
    OR2B defSlaveSMCurrentState_RNIJGOT3_inst_1 (.A(N_268), .B(
        defSlaveSMCurrentState_i_0), .Y(
        defSlaveSMCurrentState_RNIJGOT3));
    NOR2B defSlaveSMCurrentState_RNI44GI1 (.A(
        defSlaveSMCurrentState_i_0), .B(N_138), .Y(N_339));
    OR3 defSlaveSMCurrentState_RNI0ID1H (.A(N_372), .B(N_373), .C(
        N_339), .Y(N_105_i));
    NOR3C defSlaveSMNextState_i_a2_0_7 (.A(
        defSlaveSMNextState_i_a2_0_1_net_1), .B(
        defSlaveSMNextState_i_a2_0_0_net_1), .C(
        defSlaveSMNextState_i_a2_0_4_net_1), .Y(
        defSlaveSMNextState_i_a2_0_7_net_1));
    NOR3A defSlaveSMNextState_i_a2_0_6 (.A(
        defSlaveSMNextState_i_a2_0_3_net_1), .B(SDATASELInt[8]), .C(
        SDATASELInt[10]), .Y(defSlaveSMNextState_i_a2_0_6_net_1));
    VCC VCC_i (.Y(VCC));
    NOR2 defSlaveSMNextState_i_a2_0_0 (.A(SDATASELInt[9]), .B(
        SDATASELInt[13]), .Y(defSlaveSMNextState_i_a2_0_0_net_1));
    OR2 defSlaveSMCurrentState_RNISDTEF (.A(N_372), .B(N_373), .Y(
        N_261));
    NOR2 defSlaveSMNextState_i_a2_0_3 (.A(SDATASELInt[6]), .B(
        SDATASELInt[11]), .Y(defSlaveSMNextState_i_a2_0_3_net_1));
    NOR2B defSlaveSMNextState_i_a2_0 (.A(
        defSlaveSMNextState_i_a2_0_7_net_1), .B(
        defSlaveSMNextState_i_a2_0_6_net_1), .Y(N_242));
    GND GND_i (.Y(GND));
    OR2 defSlaveSMCurrentState_RNI9GQC3 (.A(N_374), .B(N_339), .Y(
        HREADY_M_iv_i_0_i_o2_0));
    OR2A defSlaveSMNextState_i_i_o2 (.A(N_242), .B(N_138), .Y(N_268));
    NOR2 defSlaveSMNextState_i_a2_0_1 (.A(SDATASELInt[12]), .B(
        SDATASELInt[15]), .Y(defSlaveSMNextState_i_a2_0_1_net_1));
    NOR2 defSlaveSMNextState_i_a2_0_4 (.A(SDATASELInt[7]), .B(
        SDATASELInt[14]), .Y(defSlaveSMNextState_i_a2_0_4_net_1));
    NOR3A defSlaveSMCurrentState_RNIMGUR2 (.A(
        defSlaveSMCurrentState_i_0), .B(m0s5DataSel), .C(N_242), .Y(
        N_373));
    
endmodule


module COREAHBLITE_MASTERSTAGE_4_1_0_32_0_1_0(
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS,
       masterAddrInProg_i_2,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE,
       HRDATA_2,
       HRDATA_1,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0,
       masterDataInProg_0,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA,
       un4_HRDATA,
       HRDATA_0_1,
       HRDATA_0_9,
       HRDATA_0_10,
       HRDATA_0_15,
       HRDATA_0_16,
       HRDATA_0_17,
       HRDATA_0_18,
       HRDATA_0_21,
       HRDATA_0_22,
       HRDATA_0_23,
       HRDATA_0_26,
       HRDATA_0_27,
       HRDATA_0_28,
       HRDATA_0_29,
       HRDATA_0_30,
       HRDATA_0_31,
       HRDATA_0_14,
       HRDATA_0_13,
       HRDATA_0_12,
       HRDATA_0_11,
       HRDATA_0_24,
       HRDATA_0_8,
       HRDATA_0_25,
       HRDATA_0_2,
       HRDATA_0_0,
       HRDATA_0_19,
       HRDATA_0_20,
       m0s5DataSel,
       masterRegAddrSel,
       defSlaveSMCurrentState_RNI5UNRI,
       CoreAHBLite_0_AHBmslave5_HREADY_i_0,
       N_63,
       N_283,
       N_284,
       N_290,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK,
       regHTRANS,
       N_259,
       N_293,
       N_292,
       N_291,
       N_153,
       FAB_CLK,
       crc_ahb_ip_MSS_0_M2F_RESET_N,
       regHWRITE,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE,
       defSlaveSMCurrentState_RNIJGOT3
    );
input  [1:1] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS;
input  [0:0] masterAddrInProg_i_2;
input  [1:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE;
input  [7:3] HRDATA_2;
input  [7:0] HRDATA_1;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0;
input  [0:0] masterDataInProg_0;
output [31:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA;
input  [31:8] un4_HRDATA;
input  HRDATA_0_1;
input  HRDATA_0_9;
input  HRDATA_0_10;
input  HRDATA_0_15;
input  HRDATA_0_16;
input  HRDATA_0_17;
input  HRDATA_0_18;
input  HRDATA_0_21;
input  HRDATA_0_22;
input  HRDATA_0_23;
input  HRDATA_0_26;
input  HRDATA_0_27;
input  HRDATA_0_28;
input  HRDATA_0_29;
input  HRDATA_0_30;
input  HRDATA_0_31;
input  HRDATA_0_14;
input  HRDATA_0_13;
input  HRDATA_0_12;
input  HRDATA_0_11;
input  HRDATA_0_24;
input  HRDATA_0_8;
input  HRDATA_0_25;
input  HRDATA_0_2;
input  HRDATA_0_0;
input  HRDATA_0_19;
input  HRDATA_0_20;
output m0s5DataSel;
output masterRegAddrSel;
output defSlaveSMCurrentState_RNI5UNRI;
input  CoreAHBLite_0_AHBmslave5_HREADY_i_0;
output N_63;
output N_283;
output N_284;
output N_290;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK;
output regHTRANS;
input  N_259;
output N_293;
output N_292;
output N_291;
output N_153;
input  FAB_CLK;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;
output regHWRITE;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE;
output defSlaveSMCurrentState_RNIJGOT3;

    wire N_371_0, N_138, d_masterRegAddrSel_0_o2_i_o2_2, 
        d_masterRegAddrSel_0_o2_i_o2_1, N_269, 
        d_masterRegAddrSel_0_i_0, N_263, d_masterRegAddrSel_0_i_o2_0_0, 
        N_285, N_264, un1_HREADY_M_pre26_1_i_i_o2_0_2, 
        \SDATASELInt[2]_net_1 , \SDATASELInt[1]_net_1 , 
        \SDATASELInt[0]_net_1 , un1_HREADY_M_pre26_1_i_i_o2_0_1, 
        \SDATASELInt[3]_net_1 , \SDATASELInt[4]_net_1 , N_375, N_280, 
        N_108, N_371, N_53, N_288, N_289, N_273, N_55, N_270, N_61, 
        N_71, N_79, \regHSIZE[0]_net_1 , \regHSIZE[1]_net_1 , 
        \regHADDR[16]_net_1 , \regHADDR[18]_net_1 , 
        \regHADDR[19]_net_1 , regHMASTLOCK_net_1, N_69, N_338, N_287, 
        \regHADDR[17]_net_1 , \regHADDR[4]_net_1 , \regHADDR[3]_net_1 , 
        \regHADDR[2]_net_1 , N_272, N_271, N_242, N_83, N_81, N_77, 
        N_75, N_73, N_67, N_65, N_59, N_57, N_374, N_372, N_105_i, 
        \SDATASELInt[6]_net_1 , \SDATASELInt[7]_net_1 , 
        \SDATASELInt[8]_net_1 , \SDATASELInt[9]_net_1 , 
        \SDATASELInt[10]_net_1 , \SDATASELInt[11]_net_1 , 
        \SDATASELInt[12]_net_1 , \SDATASELInt[13]_net_1 , 
        \SDATASELInt[14]_net_1 , \SDATASELInt[15]_net_1 , GND, VCC;
    
    NOR3 \SDATASELInt_RNO[2]  (.A(N_288), .B(N_289), .C(N_271), .Y(
        N_57));
    OA1 \SDATASELInt_RNIAEI67[5]  (.A(un4_HRDATA[25]), .B(HRDATA_0_25), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[25]));
    MX2 regHMASTLOCK_RNI5RFN (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK), .B(
        regHMASTLOCK_net_1), .S(masterRegAddrSel), .Y(N_290));
    OA1 \SDATASELInt_RNIVVJ9A[5]  (.A(HRDATA_1[6]), .B(HRDATA_2[6]), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[6]));
    OA1 \SDATASELInt_RNI48I67[5]  (.A(un4_HRDATA[22]), .B(HRDATA_0_22), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[22]));
    MX2 \regHSIZE_RNIB9FP[1]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[1]), .B(
        \regHSIZE[1]_net_1 ), .S(masterRegAddrSel), .Y(N_284));
    MX2 \regHADDR_RNIELCN[4]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2), .B(
        \regHADDR[4]_net_1 ), .S(masterRegAddrSel), .Y(N_293));
    NOR2A \SDATASELInt_RNIJ7NI1_0[5]  (.A(m0s5DataSel), .B(N_138), .Y(
        N_371));
    OA1 \SDATASELInt_RNIPQK4A[5]  (.A(HRDATA_1[5]), .B(HRDATA_2[5]), 
        .C(N_371_0), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[5])
        );
    MX2 \regHADDR_RNICJCN[2]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0), .B(
        \regHADDR[2]_net_1 ), .S(masterRegAddrSel), .Y(N_291));
    OR2A \regHADDR_RNIHNAH1[17]  (.A(N_259), .B(N_287), .Y(N_263));
    OA1 \SDATASELInt_RNI6AI67[5]  (.A(un4_HRDATA[23]), .B(HRDATA_0_23), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[23]));
    MX2 \regHADDR_RNI3B8L[18]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16), .B(
        \regHADDR[18]_net_1 ), .S(masterRegAddrSel), .Y(N_288));
    OR3 \SDATASELInt_RNI5FBP[0]  (.A(\SDATASELInt[2]_net_1 ), .B(
        \SDATASELInt[1]_net_1 ), .C(\SDATASELInt[0]_net_1 ), .Y(
        un1_HREADY_M_pre26_1_i_i_o2_0_2));
    OA1 \SDATASELInt_RNII2S77[5]  (.A(un4_HRDATA[13]), .B(HRDATA_0_13), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[13]));
    OA1 \SDATASELInt_RNI3KS77[5]  (.A(un4_HRDATA[10]), .B(HRDATA_0_10), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[10]));
    OA1 \SDATASELInt_RNI0GRC7[5]  (.A(un4_HRDATA[19]), .B(HRDATA_0_19), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[19]));
    NOR3B \SDATASELInt_RNO[14]  (.A(N_288), .B(N_289), .C(N_271), .Y(
        N_81));
    OR2 \regHADDR_RNIPT0VL[16]  (.A(d_masterRegAddrSel_0_i_o2_0_0), .B(
        N_375), .Y(N_269));
    DFN1C0 masterRegAddrSel_inst_1 (.D(N_108), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(masterRegAddrSel));
    OA1 \SDATASELInt_RNIIMI67[5]  (.A(un4_HRDATA[29]), .B(HRDATA_0_29), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[29]));
    DFN1C0 regHTRANS_inst_1 (.D(N_338), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Q(regHTRANS));
    VCC VCC_i (.Y(VCC));
    NOR3A \SDATASELInt_RNO[9]  (.A(N_289), .B(N_288), .C(N_270), .Y(
        N_71));
    OA1 \SDATASELInt_RNIUDRC7[5]  (.A(un4_HRDATA[18]), .B(HRDATA_0_18), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[18]));
    OR2 masterRegAddrSel_RNI19SB91 (.A(d_masterRegAddrSel_0_o2_i_o2_2), 
        .B(defSlaveSMCurrentState_RNI5UNRI), .Y(N_280));
    OA1 \SDATASELInt_RNINNJ9A[5]  (.A(HRDATA_1[4]), .B(HRDATA_2[4]), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[4]));
    OA1 \SDATASELInt_RNIEII67[5]  (.A(un4_HRDATA[27]), .B(HRDATA_0_27), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[27]));
    MX2 \regHADDR_RNIDKCN[3]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1), .B(
        \regHADDR[3]_net_1 ), .S(masterRegAddrSel), .Y(N_292));
    OA1 \SDATASELInt_RNI0QOG8[5]  (.A(HRDATA_0_1), .B(HRDATA_1[1]), .C(
        N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[1]));
    OR2A regHTRANS_RNO (.A(N_280), .B(regHTRANS), .Y(N_338));
    OA1 \SDATASELInt_RNIK4S77[5]  (.A(un4_HRDATA[14]), .B(HRDATA_0_14), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[14]));
    OA1 \SDATASELInt_RNICGI67[5]  (.A(un4_HRDATA[26]), .B(HRDATA_0_26), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[26]));
    OA1 \SDATASELInt_RNI8CI67[5]  (.A(un4_HRDATA[24]), .B(HRDATA_0_24), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[24]));
    MX2 \regHSIZE_RNIA8FP[0]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[0]), .B(
        \regHSIZE[0]_net_1 ), .S(masterRegAddrSel), .Y(N_283));
    NOR3A \SDATASELInt_RNO[8]  (.A(N_289), .B(N_288), .C(N_273), .Y(
        N_69));
    AO1D \SDATASELInt_RNI2KVT3[5]  (.A(N_242), .B(m0s5DataSel), .C(
        N_138), .Y(N_153));
    DFN1E0C0 \SDATASELInt[4]  (.D(N_61), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[4]_net_1 ));
    DFN1E0C0 \regHADDR[2]  (.D(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0), .CLK(FAB_CLK), 
        .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(
        \regHADDR[2]_net_1 ));
    DFN1E0C0 \SDATASELInt[15]  (.D(N_83), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[15]_net_1 ));
    NOR2 \SDATASELInt_RNO[6]  (.A(N_271), .B(N_264), .Y(N_65));
    DFN1E0C0 \SDATASELInt[14]  (.D(N_81), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[14]_net_1 ));
    MX2 \regHADDR_RNI2A8L[17]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15), .B(
        \regHADDR[17]_net_1 ), .S(masterRegAddrSel), .Y(N_287));
    DFN1E0C0 \SDATASELInt[2]  (.D(N_57), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[2]_net_1 ));
    OA1 \SDATASELInt_RNIC5OG8[5]  (.A(HRDATA_0_2), .B(HRDATA_1[2]), .C(
        N_371_0), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[2]));
    OA1 \SDATASELInt_RNIA8JR6[5]  (.A(un4_HRDATA[8]), .B(HRDATA_0_8), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[8]));
    NOR3 \SDATASELInt_RNO[3]  (.A(N_288), .B(N_289), .C(N_272), .Y(
        N_59));
    NOR3A \SDATASELInt_RNO[11]  (.A(N_289), .B(N_288), .C(N_272), .Y(
        N_75));
    NOR2A \SDATASELInt_RNI5CAQ1[5]  (.A(N_371), .B(
        masterDataInProg_0[0]), .Y(N_374));
    DFN1E0C0 \regHADDR[17]  (.D(N_269), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(
        \regHADDR[17]_net_1 ));
    GND GND_i (.Y(GND));
    OA1 \SDATASELInt_RNI34K9A[5]  (.A(HRDATA_1[7]), .B(HRDATA_2[7]), 
        .C(N_371_0), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[7])
        );
    NOR2A \SDATASELInt_RNIJ7NI1[5]  (.A(m0s5DataSel), .B(N_138), .Y(
        N_371_0));
    DFN1E0C0 \regHADDR[16]  (.D(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14), .CLK(FAB_CLK), 
        .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(
        \regHADDR[16]_net_1 ));
    OA1 \SDATASELInt_RNI7PTC7[5]  (.A(un4_HRDATA[20]), .B(HRDATA_0_20), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[20]));
    DFN1E0C0 \SDATASELInt[13]  (.D(N_79), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[13]_net_1 ));
    OA1 \SDATASELInt_RNI9RTC7[5]  (.A(un4_HRDATA[21]), .B(HRDATA_0_21), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[21]));
    DFN1E0C0 regHWRITE_inst_1 (.D(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE), .CLK(FAB_CLK), 
        .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(regHWRITE));
    OR2 \regHADDR_RNII0J62_0[16]  (.A(N_263), .B(N_285), .Y(N_273));
    DFN1E0C0 \regHSIZE[1]  (.D(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[1]), .CLK(FAB_CLK), 
        .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(
        \regHSIZE[1]_net_1 ));
    OR3B \regHADDR_RNII0J62_0[17]  (.A(N_259), .B(N_287), .C(N_285), 
        .Y(N_271));
    DFN1E0C0 regHMASTLOCK (.D(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK), .CLK(FAB_CLK), 
        .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(
        regHMASTLOCK_net_1));
    OR2A \regHADDR_RNII0J62[16]  (.A(N_285), .B(N_263), .Y(N_270));
    DFN1E0C0 \SDATASELInt[9]  (.D(N_71), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[9]_net_1 ));
    DFN1E0C0 \SDATASELInt[1]  (.D(N_55), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[1]_net_1 ));
    DFN1E0C0 \SDATASELInt[12]  (.D(N_77), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[12]_net_1 ));
    DFN1E0C0 \SDATASELInt[0]  (.D(N_53), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[0]_net_1 ));
    NOR2A d_masterRegAddrSel_0_i_a2_0 (.A(masterAddrInProg_i_2[0]), .B(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(N_375));
    OA1 \SDATASELInt_RNITMOG8[5]  (.A(HRDATA_0_0), .B(HRDATA_1[0]), .C(
        N_371_0), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[0]));
    OR2A \regHADDR_RNI80PV1[16]  (.A(N_285), .B(N_264), .Y(
        d_masterRegAddrSel_0_i_o2_0_0));
    DFN1E0C0 \SDATASELInt[5]  (.D(N_63), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(m0s5DataSel));
    OA1 \SDATASELInt_RNIPVK67[5]  (.A(un4_HRDATA[30]), .B(HRDATA_0_30), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[30]));
    OA1 \SDATASELInt_RNIO8S77[5]  (.A(un4_HRDATA[16]), .B(HRDATA_0_16), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[16]));
    OA1 \SDATASELInt_RNICAJR6[5]  (.A(un4_HRDATA[9]), .B(HRDATA_0_9), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[9]));
    NOR3B \SDATASELInt_RNO[12]  (.A(N_288), .B(N_289), .C(N_273), .Y(
        N_77));
    OR2A \regHADDR_RNI7NGA1[18]  (.A(N_288), .B(N_289), .Y(N_264));
    DFN1E0C0 \regHADDR[3]  (.D(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1), .CLK(FAB_CLK), 
        .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(
        \regHADDR[3]_net_1 ));
    OA1 \SDATASELInt_RNIM6S77[5]  (.A(un4_HRDATA[15]), .B(HRDATA_0_15), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[15]));
    OA1 \SDATASELInt_RNIG0S77[5]  (.A(un4_HRDATA[12]), .B(HRDATA_0_12), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[12]));
    DFN1E0C0 \SDATASELInt[3]  (.D(N_59), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[3]_net_1 ));
    OA1 \SDATASELInt_RNIR1L67[5]  (.A(un4_HRDATA[31]), .B(HRDATA_0_31), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[31]));
    OR2 masterRegAddrSel_RNO_0 (.A(N_263), .B(N_269), .Y(
        d_masterRegAddrSel_0_i_0));
    OR2 \SDATASELInt_RNIJ4TG[3]  (.A(\SDATASELInt[3]_net_1 ), .B(
        \SDATASELInt[4]_net_1 ), .Y(un1_HREADY_M_pre26_1_i_i_o2_0_1));
    NOR3B \SDATASELInt_RNO[15]  (.A(N_288), .B(N_289), .C(N_272), .Y(
        N_83));
    OA1 \SDATASELInt_RNIJJJ9A[5]  (.A(HRDATA_1[3]), .B(HRDATA_2[3]), 
        .C(N_371_0), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[3])
        );
    OA1 \SDATASELInt_RNI5MS77[5]  (.A(un4_HRDATA[11]), .B(HRDATA_0_11), 
        .C(N_371_0), .Y(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[11]));
    MX2 \regHADDR_RNI4C8L[19]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17), .B(
        \regHADDR[19]_net_1 ), .S(masterRegAddrSel), .Y(N_289));
    NOR3B \SDATASELInt_RNO[13]  (.A(N_288), .B(N_289), .C(N_270), .Y(
        N_79));
    DFN1E0C0 \SDATASELInt[7]  (.D(N_67), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[7]_net_1 ));
    DFN1E0C0 \regHSIZE[0]  (.D(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[0]), .CLK(FAB_CLK), 
        .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(
        \regHSIZE[0]_net_1 ));
    OR3C \regHADDR_RNII0J62[17]  (.A(N_259), .B(N_287), .C(N_285), .Y(
        N_272));
    MX2 \regHADDR_RNI198L[16]  (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14), .B(
        \regHADDR[16]_net_1 ), .S(masterRegAddrSel), .Y(N_285));
    NOR3A \SDATASELInt_RNO[10]  (.A(N_289), .B(N_288), .C(N_271), .Y(
        N_73));
    NOR3 \SDATASELInt_RNO[0]  (.A(N_288), .B(N_289), .C(N_273), .Y(
        N_53));
    NOR2 \regHADDR_RNIPN3H3[16]  (.A(N_270), .B(N_264), .Y(N_63));
    DFN1E0C0 \SDATASELInt[6]  (.D(N_65), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[6]_net_1 ));
    OA1C masterRegAddrSel_RNO (.A(defSlaveSMCurrentState_RNI5UNRI), .B(
        masterRegAddrSel), .C(d_masterRegAddrSel_0_i_0), .Y(N_108));
    DFN1E0C0 \regHADDR[19]  (.D(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17), .CLK(FAB_CLK), 
        .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(
        \regHADDR[19]_net_1 ));
    OR2 \SDATASELInt_RNIOJ8A1[0]  (.A(un1_HREADY_M_pre26_1_i_i_o2_0_2), 
        .B(un1_HREADY_M_pre26_1_i_i_o2_0_1), .Y(N_138));
    OA1 \SDATASELInt_RNIGKI67[5]  (.A(un4_HRDATA[28]), .B(HRDATA_0_28), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[28]));
    NOR2 \SDATASELInt_RNO[4]  (.A(N_273), .B(N_264), .Y(N_61));
    DFN1E0C0 \regHADDR[18]  (.D(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16), .CLK(FAB_CLK), 
        .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(
        \regHADDR[18]_net_1 ));
    OR3A masterRegAddrSel_RNI3D3H (.A(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS[1]), .B(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15), .C(
        masterRegAddrSel), .Y(d_masterRegAddrSel_0_o2_i_o2_1));
    OA1 \SDATASELInt_RNISBRC7[5]  (.A(un4_HRDATA[17]), .B(HRDATA_0_17), 
        .C(N_371), .Y(crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[17]));
    DFN1E0C0 \SDATASELInt[11]  (.D(N_75), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[11]_net_1 ));
    NOR2B \SDATASELInt_RNI6TUIC[5]  (.A(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .B(N_371), .Y(N_372));
    DFN1E0C0 \SDATASELInt[8]  (.D(N_69), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[8]_net_1 ));
    NOR2 \SDATASELInt_RNO[7]  (.A(N_272), .B(N_264), .Y(N_67));
    NOR3 \SDATASELInt_RNO[1]  (.A(N_288), .B(N_289), .C(N_270), .Y(
        N_55));
    DFN1E0C0 \regHADDR[4]  (.D(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2), .CLK(FAB_CLK), 
        .CLR(crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_280), .Q(
        \regHADDR[4]_net_1 ));
    DFN1E0C0 \SDATASELInt[10]  (.D(N_73), .CLK(FAB_CLK), .CLR(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .E(N_105_i), .Q(
        \SDATASELInt[10]_net_1 ));
    OR2 masterRegAddrSel_RNISA4GM (.A(d_masterRegAddrSel_0_o2_i_o2_1), 
        .B(N_269), .Y(d_masterRegAddrSel_0_o2_i_o2_2));
    COREAHBLITE_DEFAULTSLAVESM_default_slave_sm default_slave_sm (
        .SDATASELInt({\SDATASELInt[15]_net_1 , \SDATASELInt[14]_net_1 , 
        \SDATASELInt[13]_net_1 , \SDATASELInt[12]_net_1 , 
        \SDATASELInt[11]_net_1 , \SDATASELInt[10]_net_1 , 
        \SDATASELInt[9]_net_1 , \SDATASELInt[8]_net_1 , 
        \SDATASELInt[7]_net_1 , \SDATASELInt[6]_net_1 }), .N_372(N_372)
        , .N_374(N_374), .defSlaveSMCurrentState_RNI5UNRI(
        defSlaveSMCurrentState_RNI5UNRI), .N_242(N_242), 
        .defSlaveSMCurrentState_RNIJGOT3(
        defSlaveSMCurrentState_RNIJGOT3), .N_138(N_138), .N_105_i(
        N_105_i), .m0s5DataSel(m0s5DataSel), .FAB_CLK(FAB_CLK), 
        .crc_ahb_ip_MSS_0_M2F_RESET_N(crc_ahb_ip_MSS_0_M2F_RESET_N));
    
endmodule


module COREAHBLITE_MATRIX4X16_4_1_0_32_0_0_0(
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE,
       HRDATA_2,
       HRDATA_1,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA,
       un4_HRDATA,
       HRDATA_0_1,
       HRDATA_0_9,
       HRDATA_0_10,
       HRDATA_0_15,
       HRDATA_0_16,
       HRDATA_0_17,
       HRDATA_0_18,
       HRDATA_0_21,
       HRDATA_0_22,
       HRDATA_0_23,
       HRDATA_0_26,
       HRDATA_0_27,
       HRDATA_0_28,
       HRDATA_0_29,
       HRDATA_0_30,
       HRDATA_0_31,
       HRDATA_0_14,
       HRDATA_0_13,
       HRDATA_0_12,
       HRDATA_0_11,
       HRDATA_0_24,
       HRDATA_0_8,
       HRDATA_0_25,
       HRDATA_0_2,
       HRDATA_0_0,
       HRDATA_0_19,
       HRDATA_0_20,
       bus_wr_25,
       bus_wr_0,
       bus_wr_1,
       bus_wr_2,
       bus_wr_16,
       bus_wr_3,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA,
       defSlaveSMCurrentState_RNI5UNRI,
       CoreAHBLite_0_AHBmslave5_HREADY_i_0,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK,
       N_153,
       FAB_CLK,
       crc_ahb_ip_MSS_0_M2F_RESET_N,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE,
       N_332,
       N_333,
       N_334,
       N_335,
       N_336,
       N_337,
       N_347,
       N_348,
       N_352,
       N_353,
       N_358,
       N_360,
       N_361,
       N_364,
       N_365,
       N_366,
       N_367,
       N_350,
       N_357,
       N_356,
       N_351,
       N_349,
       N_354,
       N_362,
       N_355,
       N_363,
       un1_masterAddrInProg_6,
       N_387,
       N_408,
       N_409,
       N_5,
       N_342,
       N_341,
       N_340
    );
input  [1:1] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS;
input  [1:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE;
input  [7:3] HRDATA_2;
input  [7:0] HRDATA_1;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0;
output [31:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA;
input  [31:8] un4_HRDATA;
input  HRDATA_0_1;
input  HRDATA_0_9;
input  HRDATA_0_10;
input  HRDATA_0_15;
input  HRDATA_0_16;
input  HRDATA_0_17;
input  HRDATA_0_18;
input  HRDATA_0_21;
input  HRDATA_0_22;
input  HRDATA_0_23;
input  HRDATA_0_26;
input  HRDATA_0_27;
input  HRDATA_0_28;
input  HRDATA_0_29;
input  HRDATA_0_30;
input  HRDATA_0_31;
input  HRDATA_0_14;
input  HRDATA_0_13;
input  HRDATA_0_12;
input  HRDATA_0_11;
input  HRDATA_0_24;
input  HRDATA_0_8;
input  HRDATA_0_25;
input  HRDATA_0_2;
input  HRDATA_0_0;
input  HRDATA_0_19;
input  HRDATA_0_20;
output bus_wr_25;
output bus_wr_0;
output bus_wr_1;
output bus_wr_2;
output bus_wr_16;
output bus_wr_3;
input  [31:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA;
output defSlaveSMCurrentState_RNI5UNRI;
input  CoreAHBLite_0_AHBmslave5_HREADY_i_0;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK;
output N_153;
input  FAB_CLK;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE;
output N_332;
output N_333;
output N_334;
output N_335;
output N_336;
output N_337;
output N_347;
output N_348;
output N_352;
output N_353;
output N_358;
output N_360;
output N_361;
output N_364;
output N_365;
output N_366;
output N_367;
output N_350;
output N_357;
output N_356;
output N_351;
output N_349;
output N_354;
output N_362;
output N_355;
output N_363;
output un1_masterAddrInProg_6;
output N_387;
output N_408;
output N_409;
output N_5;
output N_342;
output N_341;
output N_340;

    wire \masterAddrInProg_i_2[0] , \masterDataInProg_0[0] , 
        m0s5DataSel, masterRegAddrSel, N_63, N_283, N_284, N_290, 
        regHTRANS, N_259, N_293, N_292, N_291, regHWRITE, 
        defSlaveSMCurrentState_RNIJGOT3, GND, VCC;
    
    COREAHBLITE_SLAVESTAGE_slavestage_5 slavestage_5 (
        .masterDataInProg_0({\masterDataInProg_0[0] }), 
        .masterAddrInProg_i_2({\masterAddrInProg_i_2[0] }), .bus_wr_25(
        bus_wr_25), .bus_wr_0(bus_wr_0), .bus_wr_1(bus_wr_1), 
        .bus_wr_2(bus_wr_2), .bus_wr_16(bus_wr_16), .bus_wr_3(bus_wr_3)
        , .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS[1]}), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[31], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[30], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[29], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[28], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[27], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[26], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[25], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[24], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[23], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[22], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[21], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[20], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[19], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[18], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[17], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[16], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[15], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[14], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[13], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[12], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[11], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[10], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[9], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[8], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[7], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[6], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[5], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[4], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[3], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[2], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[1], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[0]}), .FAB_CLK(
        FAB_CLK), .crc_ahb_ip_MSS_0_M2F_RESET_N(
        crc_ahb_ip_MSS_0_M2F_RESET_N), 
        .CoreAHBLite_0_AHBmslave5_HREADY_i_0(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .N_332(N_332), .N_333(
        N_333), .N_334(N_334), .N_335(N_335), .N_336(N_336), .N_337(
        N_337), .N_347(N_347), .N_348(N_348), .N_352(N_352), .N_353(
        N_353), .N_358(N_358), .N_360(N_360), .N_361(N_361), .N_364(
        N_364), .N_365(N_365), .N_366(N_366), .N_367(N_367), .N_350(
        N_350), .N_357(N_357), .N_356(N_356), .N_351(N_351), .N_349(
        N_349), .N_259(N_259), .regHTRANS(regHTRANS), 
        .masterRegAddrSel(masterRegAddrSel), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE), .regHWRITE(
        regHWRITE), .defSlaveSMCurrentState_RNIJGOT3(
        defSlaveSMCurrentState_RNIJGOT3), .m0s5DataSel(m0s5DataSel), 
        .N_354(N_354), .N_362(N_362), .N_355(N_355), .N_363(N_363), 
        .N_290(N_290), .N_63(N_63), .un1_masterAddrInProg_6(
        un1_masterAddrInProg_6), .N_387(N_387), .N_408(N_408), .N_283(
        N_283), .N_409(N_409), .N_284(N_284), .N_5(N_5), .N_342(N_342), 
        .N_293(N_293), .N_341(N_341), .N_292(N_292), .N_340(N_340), 
        .N_291(N_291));
    VCC VCC_i (.Y(VCC));
    COREAHBLITE_MASTERSTAGE_4_1_0_32_0_1_0 masterstage_0 (
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS[1]}), 
        .masterAddrInProg_i_2({\masterAddrInProg_i_2[0] }), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[1], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[0]}), .HRDATA_2({
        HRDATA_2[7], HRDATA_2[6], HRDATA_2[5], HRDATA_2[4], 
        HRDATA_2[3]}), .HRDATA_1({HRDATA_1[7], HRDATA_1[6], 
        HRDATA_1[5], HRDATA_1[4], HRDATA_1[3], HRDATA_1[2], 
        HRDATA_1[1], HRDATA_1[0]}), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0), 
        .masterDataInProg_0({\masterDataInProg_0[0] }), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[31], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[30], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[29], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[28], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[27], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[26], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[25], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[24], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[23], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[22], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[21], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[20], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[19], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[18], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[17], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[16], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[15], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[14], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[13], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[12], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[11], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[10], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[9], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[8], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[7], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[6], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[5], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[4], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[3], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[2], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[1], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[0]}), .un4_HRDATA({
        un4_HRDATA[31], un4_HRDATA[30], un4_HRDATA[29], un4_HRDATA[28], 
        un4_HRDATA[27], un4_HRDATA[26], un4_HRDATA[25], un4_HRDATA[24], 
        un4_HRDATA[23], un4_HRDATA[22], un4_HRDATA[21], un4_HRDATA[20], 
        un4_HRDATA[19], un4_HRDATA[18], un4_HRDATA[17], un4_HRDATA[16], 
        un4_HRDATA[15], un4_HRDATA[14], un4_HRDATA[13], un4_HRDATA[12], 
        un4_HRDATA[11], un4_HRDATA[10], un4_HRDATA[9], un4_HRDATA[8]}), 
        .HRDATA_0_1(HRDATA_0_1), .HRDATA_0_9(HRDATA_0_9), .HRDATA_0_10(
        HRDATA_0_10), .HRDATA_0_15(HRDATA_0_15), .HRDATA_0_16(
        HRDATA_0_16), .HRDATA_0_17(HRDATA_0_17), .HRDATA_0_18(
        HRDATA_0_18), .HRDATA_0_21(HRDATA_0_21), .HRDATA_0_22(
        HRDATA_0_22), .HRDATA_0_23(HRDATA_0_23), .HRDATA_0_26(
        HRDATA_0_26), .HRDATA_0_27(HRDATA_0_27), .HRDATA_0_28(
        HRDATA_0_28), .HRDATA_0_29(HRDATA_0_29), .HRDATA_0_30(
        HRDATA_0_30), .HRDATA_0_31(HRDATA_0_31), .HRDATA_0_14(
        HRDATA_0_14), .HRDATA_0_13(HRDATA_0_13), .HRDATA_0_12(
        HRDATA_0_12), .HRDATA_0_11(HRDATA_0_11), .HRDATA_0_24(
        HRDATA_0_24), .HRDATA_0_8(HRDATA_0_8), .HRDATA_0_25(
        HRDATA_0_25), .HRDATA_0_2(HRDATA_0_2), .HRDATA_0_0(HRDATA_0_0), 
        .HRDATA_0_19(HRDATA_0_19), .HRDATA_0_20(HRDATA_0_20), 
        .m0s5DataSel(m0s5DataSel), .masterRegAddrSel(masterRegAddrSel), 
        .defSlaveSMCurrentState_RNI5UNRI(
        defSlaveSMCurrentState_RNI5UNRI), 
        .CoreAHBLite_0_AHBmslave5_HREADY_i_0(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .N_63(N_63), .N_283(
        N_283), .N_284(N_284), .N_290(N_290), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK), .regHTRANS(
        regHTRANS), .N_259(N_259), .N_293(N_293), .N_292(N_292), 
        .N_291(N_291), .N_153(N_153), .FAB_CLK(FAB_CLK), 
        .crc_ahb_ip_MSS_0_M2F_RESET_N(crc_ahb_ip_MSS_0_M2F_RESET_N), 
        .regHWRITE(regHWRITE), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE), 
        .defSlaveSMCurrentState_RNIJGOT3(
        defSlaveSMCurrentState_RNIJGOT3));
    GND GND_i (.Y(GND));
    
endmodule


module CoreAHBLite_Z3(
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE,
       HRDATA_2,
       HRDATA_1,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA,
       un4_HRDATA,
       HRDATA_0_1,
       HRDATA_0_9,
       HRDATA_0_10,
       HRDATA_0_15,
       HRDATA_0_16,
       HRDATA_0_17,
       HRDATA_0_18,
       HRDATA_0_21,
       HRDATA_0_22,
       HRDATA_0_23,
       HRDATA_0_26,
       HRDATA_0_27,
       HRDATA_0_28,
       HRDATA_0_29,
       HRDATA_0_30,
       HRDATA_0_31,
       HRDATA_0_14,
       HRDATA_0_13,
       HRDATA_0_12,
       HRDATA_0_11,
       HRDATA_0_24,
       HRDATA_0_8,
       HRDATA_0_25,
       HRDATA_0_2,
       HRDATA_0_0,
       HRDATA_0_19,
       HRDATA_0_20,
       bus_wr_25,
       bus_wr_0,
       bus_wr_1,
       bus_wr_2,
       bus_wr_16,
       bus_wr_3,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA,
       defSlaveSMCurrentState_RNI5UNRI,
       CoreAHBLite_0_AHBmslave5_HREADY_i_0,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK,
       N_153,
       FAB_CLK,
       crc_ahb_ip_MSS_0_M2F_RESET_N,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE,
       N_332,
       N_333,
       N_334,
       N_335,
       N_336,
       N_337,
       N_347,
       N_348,
       N_352,
       N_353,
       N_358,
       N_360,
       N_361,
       N_364,
       N_365,
       N_366,
       N_367,
       N_350,
       N_357,
       N_356,
       N_351,
       N_349,
       N_354,
       N_362,
       N_355,
       N_363,
       un1_masterAddrInProg_6,
       N_387,
       N_408,
       N_409,
       N_5,
       N_342,
       N_341,
       N_340
    );
input  [1:1] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS;
input  [1:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE;
input  [7:3] HRDATA_2;
input  [7:0] HRDATA_1;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0;
output [31:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA;
input  [31:8] un4_HRDATA;
input  HRDATA_0_1;
input  HRDATA_0_9;
input  HRDATA_0_10;
input  HRDATA_0_15;
input  HRDATA_0_16;
input  HRDATA_0_17;
input  HRDATA_0_18;
input  HRDATA_0_21;
input  HRDATA_0_22;
input  HRDATA_0_23;
input  HRDATA_0_26;
input  HRDATA_0_27;
input  HRDATA_0_28;
input  HRDATA_0_29;
input  HRDATA_0_30;
input  HRDATA_0_31;
input  HRDATA_0_14;
input  HRDATA_0_13;
input  HRDATA_0_12;
input  HRDATA_0_11;
input  HRDATA_0_24;
input  HRDATA_0_8;
input  HRDATA_0_25;
input  HRDATA_0_2;
input  HRDATA_0_0;
input  HRDATA_0_19;
input  HRDATA_0_20;
output bus_wr_25;
output bus_wr_0;
output bus_wr_1;
output bus_wr_2;
output bus_wr_16;
output bus_wr_3;
input  [31:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA;
output defSlaveSMCurrentState_RNI5UNRI;
input  CoreAHBLite_0_AHBmslave5_HREADY_i_0;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK;
output N_153;
input  FAB_CLK;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;
input  crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE;
output N_332;
output N_333;
output N_334;
output N_335;
output N_336;
output N_337;
output N_347;
output N_348;
output N_352;
output N_353;
output N_358;
output N_360;
output N_361;
output N_364;
output N_365;
output N_366;
output N_367;
output N_350;
output N_357;
output N_356;
output N_351;
output N_349;
output N_354;
output N_362;
output N_355;
output N_363;
output un1_masterAddrInProg_6;
output N_387;
output N_408;
output N_409;
output N_5;
output N_342;
output N_341;
output N_340;

    wire GND, VCC;
    
    COREAHBLITE_MATRIX4X16_4_1_0_32_0_0_0 matrix4x16 (
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS[1]}), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[1], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[0]}), .HRDATA_2({
        HRDATA_2[7], HRDATA_2[6], HRDATA_2[5], HRDATA_2[4], 
        HRDATA_2[3]}), .HRDATA_1({HRDATA_1[7], HRDATA_1[6], 
        HRDATA_1[5], HRDATA_1[4], HRDATA_1[3], HRDATA_1[2], 
        HRDATA_1[1], HRDATA_1[0]}), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[31], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[30], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[29], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[28], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[27], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[26], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[25], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[24], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[23], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[22], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[21], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[20], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[19], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[18], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[17], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[16], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[15], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[14], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[13], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[12], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[11], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[10], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[9], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[8], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[7], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[6], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[5], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[4], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[3], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[2], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[1], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[0]}), .un4_HRDATA({
        un4_HRDATA[31], un4_HRDATA[30], un4_HRDATA[29], un4_HRDATA[28], 
        un4_HRDATA[27], un4_HRDATA[26], un4_HRDATA[25], un4_HRDATA[24], 
        un4_HRDATA[23], un4_HRDATA[22], un4_HRDATA[21], un4_HRDATA[20], 
        un4_HRDATA[19], un4_HRDATA[18], un4_HRDATA[17], un4_HRDATA[16], 
        un4_HRDATA[15], un4_HRDATA[14], un4_HRDATA[13], un4_HRDATA[12], 
        un4_HRDATA[11], un4_HRDATA[10], un4_HRDATA[9], un4_HRDATA[8]}), 
        .HRDATA_0_1(HRDATA_0_1), .HRDATA_0_9(HRDATA_0_9), .HRDATA_0_10(
        HRDATA_0_10), .HRDATA_0_15(HRDATA_0_15), .HRDATA_0_16(
        HRDATA_0_16), .HRDATA_0_17(HRDATA_0_17), .HRDATA_0_18(
        HRDATA_0_18), .HRDATA_0_21(HRDATA_0_21), .HRDATA_0_22(
        HRDATA_0_22), .HRDATA_0_23(HRDATA_0_23), .HRDATA_0_26(
        HRDATA_0_26), .HRDATA_0_27(HRDATA_0_27), .HRDATA_0_28(
        HRDATA_0_28), .HRDATA_0_29(HRDATA_0_29), .HRDATA_0_30(
        HRDATA_0_30), .HRDATA_0_31(HRDATA_0_31), .HRDATA_0_14(
        HRDATA_0_14), .HRDATA_0_13(HRDATA_0_13), .HRDATA_0_12(
        HRDATA_0_12), .HRDATA_0_11(HRDATA_0_11), .HRDATA_0_24(
        HRDATA_0_24), .HRDATA_0_8(HRDATA_0_8), .HRDATA_0_25(
        HRDATA_0_25), .HRDATA_0_2(HRDATA_0_2), .HRDATA_0_0(HRDATA_0_0), 
        .HRDATA_0_19(HRDATA_0_19), .HRDATA_0_20(HRDATA_0_20), 
        .bus_wr_25(bus_wr_25), .bus_wr_0(bus_wr_0), .bus_wr_1(bus_wr_1)
        , .bus_wr_2(bus_wr_2), .bus_wr_16(bus_wr_16), .bus_wr_3(
        bus_wr_3), .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[31], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[30], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[29], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[28], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[27], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[26], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[25], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[24], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[23], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[22], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[21], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[20], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[19], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[18], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[17], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[16], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[15], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[14], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[13], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[12], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[11], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[10], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[9], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[8], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[7], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[6], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[5], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[4], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[3], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[2], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[1], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[0]}), 
        .defSlaveSMCurrentState_RNI5UNRI(
        defSlaveSMCurrentState_RNI5UNRI), 
        .CoreAHBLite_0_AHBmslave5_HREADY_i_0(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK), .N_153(N_153), 
        .FAB_CLK(FAB_CLK), .crc_ahb_ip_MSS_0_M2F_RESET_N(
        crc_ahb_ip_MSS_0_M2F_RESET_N), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE), .N_332(N_332), 
        .N_333(N_333), .N_334(N_334), .N_335(N_335), .N_336(N_336), 
        .N_337(N_337), .N_347(N_347), .N_348(N_348), .N_352(N_352), 
        .N_353(N_353), .N_358(N_358), .N_360(N_360), .N_361(N_361), 
        .N_364(N_364), .N_365(N_365), .N_366(N_366), .N_367(N_367), 
        .N_350(N_350), .N_357(N_357), .N_356(N_356), .N_351(N_351), 
        .N_349(N_349), .N_354(N_354), .N_362(N_362), .N_355(N_355), 
        .N_363(N_363), .un1_masterAddrInProg_6(un1_masterAddrInProg_6), 
        .N_387(N_387), .N_408(N_408), .N_409(N_409), .N_5(N_5), .N_342(
        N_342), .N_341(N_341), .N_340(N_340));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    
endmodule


module host_interface(
       rev_in_type_0,
       HRDATA_2,
       HRDATA_1,
       crc_idr_out,
       HRDATA_0_20,
       HRDATA_0_15,
       HRDATA_0_31,
       HRDATA_0_2,
       HRDATA_0_17,
       HRDATA_0_0,
       HRDATA_0_28,
       HRDATA_0_29,
       HRDATA_0_26,
       HRDATA_0_11,
       HRDATA_0_12,
       HRDATA_0_16,
       HRDATA_0_30,
       HRDATA_0_14,
       HRDATA_0_19,
       HRDATA_0_13,
       HRDATA_0_27,
       HRDATA_0_25,
       HRDATA_0_24,
       HRDATA_0_8,
       HRDATA_0_9,
       HRDATA_0_10,
       HRDATA_0_1,
       HRDATA_0_18,
       HRDATA_0_21,
       HRDATA_0_22,
       HRDATA_0_23,
       state_byte,
       crc_poly_size,
       rev_in_type,
       bus_wr_0,
       bus_wr_3,
       crc_out,
       crc_poly_out,
       un4_HRDATA_9,
       un4_HRDATA_10,
       un4_HRDATA_15,
       un4_HRDATA_16,
       un4_HRDATA_17,
       un4_HRDATA_18,
       un4_HRDATA_21,
       un4_HRDATA_22,
       un4_HRDATA_23,
       un4_HRDATA_26,
       un4_HRDATA_27,
       un4_HRDATA_28,
       un4_HRDATA_29,
       un4_HRDATA_30,
       un4_HRDATA_31,
       un4_HRDATA_14,
       un4_HRDATA_13,
       un4_HRDATA_12,
       un4_HRDATA_11,
       un4_HRDATA_24,
       un4_HRDATA_8,
       un4_HRDATA_25,
       un4_HRDATA_19,
       un4_HRDATA_20,
       crc_init_out,
       bus_size,
       FAB_CLK,
       rev_out_type_0,
       crc_poly_en_0,
       crc_init_en_0,
       CoreAHBLite_0_AHBmslave5_HREADY_i_0,
       N_347,
       buffer_full,
       buffer_write_en,
       reset_pending,
       crc_ahb_ip_MSS_0_M2F_RESET_N,
       rev_out_type,
       N_350,
       reset_chain,
       crc_poly_en,
       crc_init_en,
       N_348,
       N_349,
       crc_idr_en,
       un1_masterAddrInProg_6,
       N_5,
       N_408,
       N_409,
       N_387,
       N_340,
       N_341,
       N_342
    );
output [0:0] rev_in_type_0;
output [7:3] HRDATA_2;
output [7:0] HRDATA_1;
input  [7:0] crc_idr_out;
output HRDATA_0_20;
output HRDATA_0_15;
output HRDATA_0_31;
output HRDATA_0_2;
output HRDATA_0_17;
output HRDATA_0_0;
output HRDATA_0_28;
output HRDATA_0_29;
output HRDATA_0_26;
output HRDATA_0_11;
output HRDATA_0_12;
output HRDATA_0_16;
output HRDATA_0_30;
output HRDATA_0_14;
output HRDATA_0_19;
output HRDATA_0_13;
output HRDATA_0_27;
output HRDATA_0_25;
output HRDATA_0_24;
output HRDATA_0_8;
output HRDATA_0_9;
output HRDATA_0_10;
output HRDATA_0_1;
output HRDATA_0_18;
output HRDATA_0_21;
output HRDATA_0_22;
output HRDATA_0_23;
input  [4:4] state_byte;
output [1:0] crc_poly_size;
output [1:0] rev_in_type;
input  bus_wr_0;
input  bus_wr_3;
input  [31:0] crc_out;
input  [31:0] crc_poly_out;
output un4_HRDATA_9;
output un4_HRDATA_10;
output un4_HRDATA_15;
output un4_HRDATA_16;
output un4_HRDATA_17;
output un4_HRDATA_18;
output un4_HRDATA_21;
output un4_HRDATA_22;
output un4_HRDATA_23;
output un4_HRDATA_26;
output un4_HRDATA_27;
output un4_HRDATA_28;
output un4_HRDATA_29;
output un4_HRDATA_30;
output un4_HRDATA_31;
output un4_HRDATA_14;
output un4_HRDATA_13;
output un4_HRDATA_12;
output un4_HRDATA_11;
output un4_HRDATA_24;
output un4_HRDATA_8;
output un4_HRDATA_25;
output un4_HRDATA_19;
output un4_HRDATA_20;
input  [31:0] crc_init_out;
output [1:0] bus_size;
input  FAB_CLK;
output rev_out_type_0;
output crc_poly_en_0;
output crc_init_en_0;
output CoreAHBLite_0_AHBmslave5_HREADY_i_0;
input  N_347;
input  buffer_full;
output buffer_write_en;
input  reset_pending;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;
output rev_out_type;
input  N_350;
output reset_chain;
output crc_poly_en;
output crc_init_en;
input  N_348;
input  N_349;
output crc_idr_en;
input  un1_masterAddrInProg_6;
input  N_5;
input  N_408;
input  N_409;
input  N_387;
input  N_340;
input  N_341;
input  N_342;

    wire \crc_cr_ff_RNIP7SK2[2]_net_1 , \crc_cr_ff_RNIAGJR2[4]_net_1 , 
        crc_dr_sel_0, \haddr_pp[1]_net_1 , \haddr_pp[0]_net_1 , 
        \haddr_pp[2]_net_1 , crc_init_sel_0, crc_poly_sel_0, write_en, 
        \crc_cr_ff[3]_net_1 , un3_HREADYOUT_1, \htrans_pp[1]_net_1 , 
        hselx_pp_net_1, hwrite_pp_net_1, \un11_HRDATA[20] , 
        \un11_HRDATA[15] , \un1_HRDATA[31] , \un4_HRDATA[2] , 
        crc_idr_sel, \un11_HRDATA[2] , \un11_HRDATA[17] , 
        \un4_HRDATA[6] , \un1_HRDATA[6] , \un14_HRDATA[6] , 
        \un11_HRDATA[6] , \un4_HRDATA[0] , \un11_HRDATA[0] , 
        \un11_HRDATA[28] , \un1_HRDATA[29] , \un11_HRDATA[26] , 
        \un1_HRDATA[11] , \un11_HRDATA[12] , \un11_HRDATA[16] , 
        crc_dr_sel, \un11_HRDATA[30] , \un11_HRDATA[14] , 
        \un11_HRDATA[19] , \un4_HRDATA[4] , \un1_HRDATA[4] , 
        \un14_HRDATA[4] , \un11_HRDATA[4] , \un1_HRDATA[13] , 
        \un1_HRDATA[7] , \un4_HRDATA[7] , \un14_HRDATA[7] , 
        \un11_HRDATA[7] , \un1_HRDATA[27] , \un11_HRDATA[25] , 
        \un11_HRDATA[24] , \un1_HRDATA[8] , \un1_HRDATA[9] , 
        \un11_HRDATA[10] , \un4_HRDATA[3] , \un1_HRDATA[3] , 
        \un14_HRDATA[3] , \un11_HRDATA[3] , crc_cr_sel, \HRDATA_0[5] , 
        \un11_HRDATA[5] , \un4_HRDATA[5] , \un4_HRDATA[1] , 
        \un11_HRDATA[1] , \un1_HRDATA[18] , \un11_HRDATA[21] , 
        \un11_HRDATA[22] , \un1_HRDATA[23] , un3_HREADYOUT, 
        crc_init_sel, un4_HREADYOUT, un2_HREADYOUT, crc_poly_sel, 
        N_364, crc_cr_en, hselx_pp5, \crc_cr_ff_RNO[1]_net_1 , N_367, 
        N_365, N_363, N_366, \crc_cr_ff_RNO[0]_net_1 , 
        \crc_cr_ff_RNO[3]_net_1 , hselx_pp_RNO_net_1, N_362, GND, VCC;
    
    DFN1 hselx_pp (.D(hselx_pp_RNO_net_1), .CLK(FAB_CLK), .Q(
        hselx_pp_net_1));
    NOR2B hwrite_pp_RNI4SA52_4 (.A(write_en), .B(crc_idr_sel), .Y(
        crc_idr_en));
    NOR2B \haddr_pp_RNIQK1M1[0]  (.A(crc_init_out[18]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_18));
    NOR3B \haddr_pp_RNISEFF1_0[0]  (.A(\haddr_pp[2]_net_1 ), .B(
        \haddr_pp[0]_net_1 ), .C(\haddr_pp[1]_net_1 ), .Y(crc_poly_sel)
        );
    OR3 \haddr_pp_RNI3PHD5[0]  (.A(\un4_HRDATA[6] ), .B(
        \un1_HRDATA[6] ), .C(\un14_HRDATA[6] ), .Y(HRDATA_2[6]));
    AO1 \crc_cr_ff_0_0_RNIVLI85[2]  (.A(crc_cr_sel), .B(
        rev_in_type_0[0]), .C(\HRDATA_0[5] ), .Y(HRDATA_2[5]));
    NOR3A \haddr_pp_RNISEFF1_1[0]  (.A(\haddr_pp[0]_net_1 ), .B(
        \haddr_pp[1]_net_1 ), .C(\haddr_pp[2]_net_1 ), .Y(crc_idr_sel));
    NOR2B \haddr_pp_RNIIC5K1[0]  (.A(crc_poly_out[1]), .B(
        crc_poly_sel_0), .Y(\un11_HRDATA[1] ));
    NOR2B \haddr_pp_RNI4P1Q1[0]  (.A(crc_poly_out[12]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[12] ));
    DFN1 \crc_cr_ff[2]  (.D(\crc_cr_ff_RNIP7SK2[2]_net_1 ), .CLK(
        FAB_CLK), .Q(rev_in_type[0]));
    AO1 \haddr_pp_RNI1NA93[0]  (.A(crc_idr_out[2]), .B(crc_idr_sel), 
        .C(\un11_HRDATA[2] ), .Y(HRDATA_0_2));
    NOR2B \haddr_pp_RNIJD5K1[0]  (.A(crc_poly_out[2]), .B(
        crc_poly_sel_0), .Y(\un11_HRDATA[2] ));
    NOR2B \haddr_pp_RNI6R1Q1[0]  (.A(crc_poly_out[14]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[14] ));
    NOR2B \haddr_pp_RNI9PVL1[0]  (.A(crc_init_out[8]), .B(crc_init_sel)
        , .Y(un4_HRDATA_8));
    NOR2B \haddr_pp_RNIKG3M1[0]  (.A(crc_init_out[30]), .B(
        crc_init_sel), .Y(un4_HRDATA_30));
    AO1 \haddr_pp_RNITGOT3[0]  (.A(crc_poly_out[23]), .B(
        crc_poly_sel_0), .C(\un1_HRDATA[23] ), .Y(HRDATA_0_23));
    AO1 \haddr_pp_RNI3PA93[0]  (.A(crc_idr_out[3]), .B(crc_idr_sel), 
        .C(\un11_HRDATA[3] ), .Y(HRDATA_1[3]));
    NOR2B hwrite_pp_RNI4SA52_1 (.A(write_en), .B(crc_poly_sel), .Y(
        crc_poly_en));
    NOR2B \haddr_pp_RNIAQVL1[0]  (.A(crc_init_out[9]), .B(crc_init_sel)
        , .Y(un4_HRDATA_9));
    NOR2B \haddr_pp_RNI5H152[0]  (.A(crc_out[13]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[13] ));
    NOR3 \haddr_pp_RNISEFF1_5[0]  (.A(\haddr_pp[1]_net_1 ), .B(
        \haddr_pp[0]_net_1 ), .C(\haddr_pp[2]_net_1 ), .Y(crc_dr_sel_0)
        );
    NOR2B \haddr_pp_RNI7S1Q1[0]  (.A(crc_poly_out[15]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[15] ));
    NOR2B \haddr_pp_RNIOI5K1[0]  (.A(crc_poly_out[7]), .B(crc_poly_sel)
        , .Y(\un11_HRDATA[7] ));
    DFN1 \crc_cr_ff[4]  (.D(\crc_cr_ff_RNIAGJR2[4]_net_1 ), .CLK(
        FAB_CLK), .Q(rev_out_type));
    NOR2B \crc_cr_ff_RNI5CRO1[1]  (.A(crc_poly_size[1]), .B(crc_cr_sel)
        , .Y(\un14_HRDATA[4] ));
    DFN1E1 \hsize_pp[0]  (.D(N_408), .CLK(FAB_CLK), .E(hselx_pp5), .Q(
        bus_size[0]));
    NOR2B \haddr_pp_RNI1HVL1[0]  (.A(crc_init_out[0]), .B(crc_init_sel)
        , .Y(\un4_HRDATA[0] ));
    NOR2B \haddr_pp_RNI2IVL1[0]  (.A(crc_init_out[1]), .B(crc_init_sel)
        , .Y(\un4_HRDATA[1] ));
    NOR2B \haddr_pp_RNIQL2M1[0]  (.A(crc_init_out[27]), .B(
        crc_init_sel), .Y(un4_HRDATA_27));
    NOR2B \haddr_pp_RNILJMU1_1[0]  (.A(crc_out[3]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[3] ));
    AO1 \haddr_pp_RNI13444[0]  (.A(crc_out[20]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[20] ), .Y(HRDATA_0_20));
    NOR2B hwrite_pp_RNI4SA52 (.A(write_en), .B(crc_init_sel_0), .Y(
        crc_init_en));
    NOR2B \haddr_pp_RNIOI1M1[0]  (.A(crc_init_out[16]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_16));
    NOR2B hwrite_pp_RNI4SA52_3 (.A(write_en), .B(crc_dr_sel), .Y(
        buffer_write_en));
    OR3 hwrite_pp_RNIJL70B (.A(un4_HREADYOUT), .B(un3_HREADYOUT), .C(
        un2_HREADYOUT), .Y(CoreAHBLite_0_AHBmslave5_HREADY_i_0));
    NOR2B \haddr_pp_RNIRL1M1[0]  (.A(crc_init_out[19]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_19));
    DFN1E1 \hsize_pp[1]  (.D(N_409), .CLK(FAB_CLK), .E(hselx_pp5), .Q(
        bus_size[1]));
    NOR2B \haddr_pp_RNIKE5K1[0]  (.A(crc_poly_out[3]), .B(
        crc_poly_sel_0), .Y(\un11_HRDATA[3] ));
    NOR2B \haddr_pp_RNI9U1Q1[0]  (.A(crc_poly_out[17]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[17] ));
    DFN1E1 \haddr_pp[0]  (.D(N_340), .CLK(FAB_CLK), .E(hselx_pp5), .Q(
        \haddr_pp[0]_net_1 ));
    GND GND_i (.Y(GND));
    NOR2B hselx_pp_RNO (.A(N_362), .B(crc_ahb_ip_MSS_0_M2F_RESET_N), 
        .Y(hselx_pp_RNO_net_1));
    NOR2B \haddr_pp_RNISN2M1[0]  (.A(crc_init_out[29]), .B(
        crc_init_sel), .Y(un4_HRDATA_29));
    AO1 \haddr_pp_RNIII244[0]  (.A(crc_out[19]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[19] ), .Y(HRDATA_0_19));
    NOR2B \haddr_pp_RNI7NVL1[0]  (.A(crc_init_out[6]), .B(crc_init_sel)
        , .Y(\un4_HRDATA[6] ));
    NOR2B \haddr_pp_RNILJMU1_4[0]  (.A(crc_out[8]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[8] ));
    DFN1 \crc_cr_ff_0_0[4]  (.D(\crc_cr_ff_RNIAGJR2[4]_net_1 ), .CLK(
        FAB_CLK), .Q(rev_out_type_0));
    NOR3B \haddr_pp_RNISEFF1[0]  (.A(\haddr_pp[2]_net_1 ), .B(
        \haddr_pp[0]_net_1 ), .C(\haddr_pp[1]_net_1 ), .Y(
        crc_poly_sel_0));
    NOR2B \haddr_pp_RNIRHR82[0]  (.A(crc_cr_en), .B(bus_wr_0), .Y(
        reset_chain));
    NOR2B \haddr_pp_RNIOJ2M1[0]  (.A(crc_init_out[25]), .B(
        crc_init_sel), .Y(un4_HRDATA_25));
    NOR2B \haddr_pp_RNI2N1Q1[0]  (.A(crc_poly_out[10]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[10] ));
    NOR2B \haddr_pp_RNILF1M1[0]  (.A(crc_init_out[13]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_13));
    MX2 \crc_cr_ff_RNIMOUO2[4]  (.A(rev_out_type), .B(N_350), .S(
        crc_cr_en), .Y(N_367));
    AO1 \haddr_pp_RNIV04V3[0]  (.A(crc_poly_out[11]), .B(
        crc_poly_sel_0), .C(\un1_HRDATA[11] ), .Y(HRDATA_0_11));
    NOR2B \haddr_pp_RNINKL32[0]  (.A(crc_out[29]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[29] ));
    NOR2B \haddr_pp_RNIKE1M1[0]  (.A(crc_init_out[12]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_12));
    AO1 \haddr_pp_RNIUHOT3[0]  (.A(crc_out[24]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[24] ), .Y(HRDATA_0_24));
    NOR3B hwrite_pp_RNI8DRL_0 (.A(\htrans_pp[1]_net_1 ), .B(
        hselx_pp_net_1), .C(hwrite_pp_net_1), .Y(un3_HREADYOUT_1));
    NOR2B \haddr_pp_RNIECM32[0]  (.A(crc_out[31]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[31] ));
    AO1 \haddr_pp_RNIO6MK3[0]  (.A(crc_out[2]), .B(crc_dr_sel_0), .C(
        \un4_HRDATA[2] ), .Y(HRDATA_1[2]));
    AO1 \haddr_pp_RNII7QT3[0]  (.A(crc_out[30]), .B(crc_dr_sel), .C(
        \un11_HRDATA[30] ), .Y(HRDATA_0_30));
    AO1 \haddr_pp_RNI0KOT3[0]  (.A(crc_out[26]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[26] ), .Y(HRDATA_0_26));
    AO1 \haddr_pp_RNIBC3V3[0]  (.A(crc_out[14]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[14] ), .Y(HRDATA_0_14));
    NOR2B \haddr_pp_RNINH1M1[0]  (.A(crc_init_out[15]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_15));
    AO1 \haddr_pp_RNIHH244[0]  (.A(crc_poly_out[18]), .B(
        crc_poly_sel_0), .C(\un1_HRDATA[18] ), .Y(HRDATA_0_18));
    VCC VCC_i (.Y(VCC));
    NOR2B \haddr_pp_RNIS8252[0]  (.A(crc_out[11]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[11] ));
    AO1 \haddr_pp_RNIETMK3[0]  (.A(crc_out[1]), .B(crc_dr_sel_0), .C(
        \un4_HRDATA[1] ), .Y(HRDATA_1[1]));
    NOR2B \haddr_pp_RNILJMU1_3[0]  (.A(crc_out[9]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[9] ));
    NOR2B \haddr_pp_RNIIC1M1[0]  (.A(crc_init_out[10]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_10));
    NOR2B \haddr_pp_RNINI2M1[0]  (.A(crc_init_out[24]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_24));
    NOR2B \haddr_pp_RNILJMU1_0[0]  (.A(crc_out[4]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[4] ));
    AO1 \haddr_pp_RNI24444[0]  (.A(crc_out[21]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[21] ), .Y(HRDATA_0_21));
    AO1 \haddr_pp_RNIAB3V3[0]  (.A(crc_poly_out[13]), .B(
        crc_poly_sel_0), .C(\un1_HRDATA[13] ), .Y(HRDATA_0_13));
    DFN1E1 \haddr_pp[1]  (.D(N_341), .CLK(FAB_CLK), .E(hselx_pp5), .Q(
        \haddr_pp[1]_net_1 ));
    NOR2B \haddr_pp_RNINH5K1[0]  (.A(crc_poly_out[6]), .B(
        crc_poly_sel_0), .Y(\un11_HRDATA[6] ));
    NOR2B \haddr_pp_RNINKL32_0[0]  (.A(crc_out[27]), .B(crc_dr_sel), 
        .Y(\un1_HRDATA[27] ));
    MX2A hselx_pp_RNO_0 (.A(un1_masterAddrInProg_6), .B(hselx_pp_net_1)
        , .S(CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(N_362));
    OR3 \crc_cr_ff_RNIVKHD5[1]  (.A(\un4_HRDATA[4] ), .B(
        \un1_HRDATA[4] ), .C(\un14_HRDATA[4] ), .Y(HRDATA_2[4]));
    AO1 \haddr_pp_RNITIA93[0]  (.A(crc_idr_out[0]), .B(crc_idr_sel), 
        .C(\un11_HRDATA[0] ), .Y(HRDATA_0_0));
    AO1 \haddr_pp_RNIDE3V3[0]  (.A(crc_out[16]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[16] ), .Y(HRDATA_0_16));
    NOR2B hwrite_pp_RNINT8D2 (.A(reset_pending), .B(crc_init_en_0), .Y(
        un4_HREADYOUT));
    NOR2B \haddr_pp_RNI8U2Q1[0]  (.A(crc_poly_out[25]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[25] ));
    NOR2B hwrite_pp_RNI4SA52_0 (.A(write_en), .B(crc_init_sel_0), .Y(
        crc_init_en_0));
    NOR2B \crc_cr_ff_RNI8FRO1[4]  (.A(crc_cr_sel), .B(rev_out_type), 
        .Y(\un14_HRDATA[7] ));
    AO1 \haddr_pp_RNI5RA93[0]  (.A(crc_idr_out[4]), .B(crc_idr_sel), 
        .C(\un11_HRDATA[4] ), .Y(HRDATA_1[4]));
    NOR2B \haddr_pp_RNIPK2M1[0]  (.A(crc_init_out[26]), .B(
        crc_init_sel), .Y(un4_HRDATA_26));
    NOR2B \crc_cr_ff_RNI4BRO1[0]  (.A(crc_poly_size[0]), .B(crc_cr_sel)
        , .Y(\un14_HRDATA[3] ));
    NOR2B \haddr_pp_RNI5R2Q1[0]  (.A(crc_poly_out[22]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[22] ));
    NOR2B \haddr_pp_RNI4Q2Q1[0]  (.A(crc_poly_out[21]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[21] ));
    NOR2B \haddr_pp_RNILJMU1[0]  (.A(crc_out[6]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[6] ));
    NOR3A \haddr_pp_RNISEFF1_4[0]  (.A(\haddr_pp[1]_net_1 ), .B(
        \haddr_pp[0]_net_1 ), .C(\haddr_pp[2]_net_1 ), .Y(crc_cr_sel));
    AO1 \haddr_pp_RNISFOT3[0]  (.A(crc_out[22]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[22] ), .Y(HRDATA_0_22));
    AO1 \haddr_pp_RNI9A3V3[0]  (.A(crc_out[12]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[12] ), .Y(HRDATA_0_12));
    MX2 \crc_cr_ff_RNI5G7I2[2]  (.A(rev_in_type[0]), .B(N_348), .S(
        crc_cr_en), .Y(N_365));
    NOR2B \haddr_pp_RNIHB5K1[0]  (.A(crc_poly_out[0]), .B(
        crc_poly_sel_0), .Y(\un11_HRDATA[0] ));
    NOR2A hwrite_pp_RNI7DS2B (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .Y(hselx_pp5));
    NOR2B \haddr_pp_RNI5LVL1[0]  (.A(crc_init_out[4]), .B(crc_init_sel)
        , .Y(\un4_HRDATA[4] ));
    AO1 \haddr_pp_RNIR9MK3[0]  (.A(crc_out[5]), .B(crc_dr_sel), .C(
        \un4_HRDATA[5] ), .Y(\HRDATA_0[5] ));
    NOR2B \haddr_pp_RNIPJ1M1[0]  (.A(crc_init_out[17]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_17));
    NOR2B \haddr_pp_RNI9V2Q1[0]  (.A(crc_poly_out[26]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[26] ));
    NOR3 \haddr_pp_RNISEFF1_6[0]  (.A(\haddr_pp[1]_net_1 ), .B(
        \haddr_pp[0]_net_1 ), .C(\haddr_pp[2]_net_1 ), .Y(crc_dr_sel));
    DFN1E1 \htrans_pp[1]  (.D(N_387), .CLK(FAB_CLK), .E(hselx_pp5), .Q(
        \htrans_pp[1]_net_1 ));
    AO1 \haddr_pp_RNI7TA93[0]  (.A(crc_idr_out[5]), .B(crc_idr_sel), 
        .C(\un11_HRDATA[5] ), .Y(HRDATA_1[5]));
    NOR2B \haddr_pp_RNI4KVL1[0]  (.A(crc_init_out[3]), .B(crc_init_sel)
        , .Y(\un4_HRDATA[3] ));
    NOR2B hwrite_pp_RNIOVG56 (.A(buffer_full), .B(buffer_write_en), .Y(
        un2_HREADYOUT));
    MX2 \crc_cr_ff_RNO_0[1]  (.A(crc_poly_size[1]), .B(N_347), .S(
        crc_cr_en), .Y(N_364));
    AO1 \haddr_pp_RNIE7SI3[0]  (.A(crc_poly_out[8]), .B(crc_poly_sel_0)
        , .C(\un1_HRDATA[8] ), .Y(HRDATA_0_8));
    NOR2B \haddr_pp_RNILJMU1_2[0]  (.A(crc_out[7]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[7] ));
    NOR3A \haddr_pp_RNISEFF1_3[0]  (.A(\haddr_pp[2]_net_1 ), .B(
        \haddr_pp[0]_net_1 ), .C(\haddr_pp[1]_net_1 ), .Y(crc_init_sel)
        );
    NOR2B \haddr_pp_RNIB13Q1[0]  (.A(crc_poly_out[28]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[28] ));
    DFN1E1 \haddr_pp[2]  (.D(N_342), .CLK(FAB_CLK), .E(hselx_pp5), .Q(
        \haddr_pp[2]_net_1 ));
    MX2 \crc_cr_ff_RNO_0[0]  (.A(crc_poly_size[0]), .B(bus_wr_3), .S(
        crc_cr_en), .Y(N_363));
    NOR2B \haddr_pp_RNI7I0A2[0]  (.A(crc_out[18]), .B(crc_dr_sel), .Y(
        \un1_HRDATA[18] ));
    NOR2B \haddr_pp_RNI7ERO1[0]  (.A(crc_cr_sel), .B(rev_in_type[1]), 
        .Y(\un14_HRDATA[6] ));
    NOR3B hwrite_pp_RNI4ODD2 (.A(un3_HREADYOUT_1), .B(crc_dr_sel), .C(
        state_byte[4]), .Y(un3_HREADYOUT));
    AO1 \haddr_pp_RNI3NOT3[0]  (.A(crc_poly_out[29]), .B(
        crc_poly_sel_0), .C(\un1_HRDATA[29] ), .Y(HRDATA_0_29));
    DFN1 \crc_cr_ff[1]  (.D(\crc_cr_ff_RNO[1]_net_1 ), .CLK(FAB_CLK), 
        .Q(crc_poly_size[1]));
    AO1 \haddr_pp_RNICD3V3[0]  (.A(crc_out[15]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[15] ), .Y(HRDATA_0_15));
    NOR2B \crc_cr_ff_RNIP7SK2[2]  (.A(N_365), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(
        \crc_cr_ff_RNIP7SK2[2]_net_1 ));
    NOR2B \haddr_pp_RNILH3M1[0]  (.A(crc_init_out[31]), .B(
        crc_init_sel), .Y(un4_HRDATA_31));
    DFN1 \crc_cr_ff[3]  (.D(\crc_cr_ff_RNO[3]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_cr_ff[3]_net_1 ));
    NOR2B \haddr_pp_RNI7T2Q1[0]  (.A(crc_poly_out[24]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[24] ));
    OR3 \crc_cr_ff_RNI5RHD5[4]  (.A(\un1_HRDATA[7] ), .B(
        \un4_HRDATA[7] ), .C(\un14_HRDATA[7] ), .Y(HRDATA_2[7]));
    NOR2B \haddr_pp_RNI8T1Q1[0]  (.A(crc_poly_out[16]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[16] ));
    NOR2B \haddr_pp_RNIKF2M1[0]  (.A(crc_init_out[21]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_21));
    NOR2B \haddr_pp_RNIB02Q1[0]  (.A(crc_poly_out[19]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[19] ));
    DFN1 \crc_cr_ff[0]  (.D(\crc_cr_ff_RNO[0]_net_1 ), .CLK(FAB_CLK), 
        .Q(crc_poly_size[0]));
    NOR2B \haddr_pp_RNI6MVL1[0]  (.A(crc_init_out[5]), .B(crc_init_sel)
        , .Y(\un4_HRDATA[5] ));
    AO1 \haddr_pp_RNIJ8QT3[0]  (.A(crc_poly_out[31]), .B(
        crc_poly_sel_0), .C(\un1_HRDATA[31] ), .Y(HRDATA_0_31));
    NOR2B hwrite_pp_RNI4SA52_2 (.A(write_en), .B(crc_poly_sel_0), .Y(
        crc_poly_en_0));
    NOR2B \haddr_pp_RNIRM2M1[0]  (.A(crc_init_out[28]), .B(
        crc_init_sel), .Y(un4_HRDATA_28));
    NOR2B \crc_cr_ff_RNO[3]  (.A(N_366), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_cr_ff_RNO[3]_net_1 ));
    AO1 \haddr_pp_RNIB1B93[0]  (.A(crc_idr_out[7]), .B(crc_idr_sel), 
        .C(\un11_HRDATA[7] ), .Y(HRDATA_1[7]));
    DFN1 \crc_cr_ff_0_0[2]  (.D(\crc_cr_ff_RNIP7SK2[2]_net_1 ), .CLK(
        FAB_CLK), .Q(rev_in_type_0[0]));
    NOR2B \haddr_pp_RNIMG1M1[0]  (.A(crc_init_out[14]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_14));
    NOR2B \haddr_pp_RNI8OVL1[0]  (.A(crc_init_out[7]), .B(crc_init_sel)
        , .Y(\un4_HRDATA[7] ));
    NOR2B \haddr_pp_RNI4SA52[0]  (.A(write_en), .B(crc_cr_sel), .Y(
        crc_cr_en));
    NOR2B \haddr_pp_RNIJE2M1[0]  (.A(crc_init_out[20]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_20));
    DFN1E1 hwrite_pp (.D(N_5), .CLK(FAB_CLK), .E(hselx_pp5), .Q(
        hwrite_pp_net_1));
    AO1 \haddr_pp_RNI2MOT3[0]  (.A(crc_out[28]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[28] ), .Y(HRDATA_0_28));
    NOR3A \haddr_pp_RNISEFF1_2[0]  (.A(\haddr_pp[2]_net_1 ), .B(
        \haddr_pp[0]_net_1 ), .C(\haddr_pp[1]_net_1 ), .Y(
        crc_init_sel_0));
    OR3 \crc_cr_ff_RNITIHD5[0]  (.A(\un4_HRDATA[3] ), .B(
        \un1_HRDATA[3] ), .C(\un14_HRDATA[3] ), .Y(HRDATA_2[3]));
    NOR2B \haddr_pp_RNI3JVL1[0]  (.A(crc_init_out[2]), .B(crc_init_sel)
        , .Y(\un4_HRDATA[2] ));
    NOR2B \crc_cr_ff_RNO[1]  (.A(N_364), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_cr_ff_RNO[1]_net_1 ));
    NOR2B \haddr_pp_RNI3P2Q1[0]  (.A(crc_poly_out[20]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[20] ));
    CLKINT \crc_cr_ff_RNIBVB9[3]  (.A(\crc_cr_ff[3]_net_1 ), .Y(
        rev_in_type[1]));
    AO1 \haddr_pp_RNIVIOT3[0]  (.A(crc_out[25]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[25] ), .Y(HRDATA_0_25));
    NOR2B \haddr_pp_RNIMH2M1[0]  (.A(crc_init_out[23]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_23));
    AO1 \haddr_pp_RNIUV3V3[0]  (.A(crc_out[10]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[10] ), .Y(HRDATA_0_10));
    NOR2B \haddr_pp_RNILF5K1[0]  (.A(crc_poly_out[4]), .B(
        crc_poly_sel_0), .Y(\un11_HRDATA[4] ));
    NOR2B \crc_cr_ff_RNO[0]  (.A(N_363), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_cr_ff_RNO[0]_net_1 ));
    AO1 \haddr_pp_RNI9VA93[0]  (.A(crc_idr_out[6]), .B(crc_idr_sel), 
        .C(\un11_HRDATA[6] ), .Y(HRDATA_1[6]));
    NOR2B \crc_cr_ff_RNIAGJR2[4]  (.A(N_367), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(
        \crc_cr_ff_RNIAGJR2[4]_net_1 ));
    AO1 \haddr_pp_RNIVKA93[0]  (.A(crc_idr_out[1]), .B(crc_idr_sel), 
        .C(\un11_HRDATA[1] ), .Y(HRDATA_0_1));
    AO1 \haddr_pp_RNI1LOT3[0]  (.A(crc_poly_out[27]), .B(
        crc_poly_sel_0), .C(\un1_HRDATA[27] ), .Y(HRDATA_0_27));
    MX2 \crc_cr_ff_RNO_0[3]  (.A(rev_in_type[1]), .B(N_349), .S(
        crc_cr_en), .Y(N_366));
    AO1 \haddr_pp_RNIF8SI3[0]  (.A(crc_poly_out[9]), .B(crc_poly_sel_0)
        , .C(\un1_HRDATA[9] ), .Y(HRDATA_0_9));
    NOR3C hwrite_pp_RNI8DRL (.A(\htrans_pp[1]_net_1 ), .B(
        hselx_pp_net_1), .C(hwrite_pp_net_1), .Y(write_en));
    NOR2B \haddr_pp_RNIJD1M1[0]  (.A(crc_init_out[11]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_11));
    NOR2B \haddr_pp_RNI4R3Q1[0]  (.A(crc_poly_out[30]), .B(
        crc_poly_sel), .Y(\un11_HRDATA[30] ));
    NOR2B \haddr_pp_RNILG2M1[0]  (.A(crc_init_out[22]), .B(
        crc_init_sel_0), .Y(un4_HRDATA_22));
    NOR2B \haddr_pp_RNINKL32_1[0]  (.A(crc_out[23]), .B(crc_dr_sel), 
        .Y(\un1_HRDATA[23] ));
    NOR2B \haddr_pp_RNIMG5K1[0]  (.A(crc_poly_out[5]), .B(
        crc_poly_sel_0), .Y(\un11_HRDATA[5] ));
    AO1 \haddr_pp_RNIDSMK3[0]  (.A(crc_out[0]), .B(crc_dr_sel_0), .C(
        \un4_HRDATA[0] ), .Y(HRDATA_1[0]));
    AO1 \haddr_pp_RNIGG244[0]  (.A(crc_out[17]), .B(crc_dr_sel_0), .C(
        \un11_HRDATA[17] ), .Y(HRDATA_0_17));
    
endmodule


module crc_control_unit(
       state_byte_0,
       size_in,
       state_byte_3,
       state_byte_i,
       FAB_CLK,
       byte_en_0,
       buffer_en_0,
       buffer_write_en,
       buffer_full,
       reset_pending,
       reset_chain,
       N_294,
       crc_ahb_ip_MSS_0_M2F_RESET_N,
       N_128,
       byte_en,
       N_56,
       bypass_byte0,
       buffer_en,
       N_118_1
    );
output [4:4] state_byte_0;
input  [1:0] size_in;
output state_byte_3;
output [0:0] state_byte_i;
input  FAB_CLK;
output byte_en_0;
output buffer_en_0;
input  buffer_write_en;
output buffer_full;
output reset_pending;
input  reset_chain;
output N_294;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;
output N_128;
output byte_en;
output N_56;
output bypass_byte0;
output buffer_en;
output N_118_1;

    wire \state_byte_nss[4] , N_54, \state_full[1]_net_1 , N_118, 
        \state_reset_ns_i_a2_i_0_2[1] , \state_reset_ns_i_a2_i_0_0[1] , 
        N_135, \state_reset_RNO_4[1]_net_1 , N_165, N_1006_tz, 
        \state_reset_RNO_6[1]_net_1 , \state_reset_ns_i_a2_i_0_3[0] , 
        N_110, \state_reset[1]_net_1 , \state_reset_ns_i_a2_i_0_2[0] , 
        N_148, N_151, \state_reset_ns_i_a2_i_0_0[0] , N_153, 
        \state_full_ns_i_i_0_1[0]_net_1 , N_55, 
        \state_full_ns_i_i_0_0[0]_net_1 , \state_full[0]_net_1 , 
        \state_reset_ns_i_a2_0_0_0[4] , \state_reset[3]_net_1 , 
        \state_reset[4]_net_1 , \state_reset_ns_i_a2_i_0_a7_0_0[3] , 
        N_70, \state_reset_ns_i_a2_i_0_o2_1_0[3] , N_434, N_173, 
        \state_byte_ns_i_0_0_2[0] , \state_byte_ns_i_0_0_0[0] , 
        \state_byte_ns[2] , \state_byte[2]_net_1 , 
        \state_byte_ns_0_0_0_0[4] , N_134, 
        \state_reset_ns_i_a2_i_0_a7_0[0] , 
        state_reset_ns_i_a2_i_0_125_tz_0, N_438, 
        \state_reset_ns_i_a2_i_0_a7_7_0[1] , 
        \state_reset_ns_i_a2_i_0_a7_2_0[0] , 
        \state_reset_ns_i_a2_i_0_a7_4_0[0] , 
        clear_crc_init_sel_i_0_a7_0, \state_reset_ns_i_a2_0_0_o2_0[2] , 
        N_133, N_435, N_102, N_430, N_167, N_155, 
        \state_byte[3]_net_1 , N_154, N_95, N_146, N_137, N_124, N_177, 
        N_123, \state_reset_ns_i_a2_i_0_a7_8_0[1] , 
        \state_reset_ns_i_a2_i_0_a7_2_0[1] , N_1004_tz, N_169, 
        \state_byte[1]_net_1 , \state_full_nss[0] , 
        \state_full_nss[1] , N_122, \state_reset_nss[0] , N_150, 
        \state_reset_nss[1] , \state_reset_nss[2] , N_129, 
        \state_reset_nss[3] , N_4, \state_reset_nss[4] , 
        \state_byte_nss[0] , \state_byte_ns[1] , \state_byte_nss[1] , 
        \state_byte_nss[2] , \state_byte_nss[3] , N_125, 
        \state_reset[2]_net_1 , N_160, N_111, N_174, N_176, N_157, 
        N_159, N_166, N_431, N_64, GND, VCC;
    
    NOR2A \state_reset_RNO_7[1]  (.A(N_165), .B(state_byte_3), .Y(
        N_160));
    NOR2B \state_reset_RNO_14[1]  (.A(\state_byte[3]_net_1 ), .B(
        size_in[0]), .Y(\state_reset_ns_i_a2_i_0_a7_7_0[1] ));
    OR2A \state_reset_i_RNIFJPE[0]  (.A(\state_full[1]_net_1 ), .B(
        reset_pending), .Y(\state_reset_ns_i_a2_0_0_o2_0[2] ));
    NOR3C \state_full_ns_0_i_i_a7_0[1]  (.A(buffer_write_en), .B(
        \state_full[0]_net_1 ), .C(N_54), .Y(N_123));
    NOR2B \state_reset_RNO_1[3]  (.A(N_70), .B(buffer_write_en), .Y(
        \state_reset_ns_i_a2_i_0_a7_0_0[3] ));
    OR2 \state_byte_RNIAIFEA[4]  (.A(N_124), .B(N_125), .Y(N_56));
    AO1A \state_byte_i_RNO_1[0]  (.A(buffer_write_en), .B(
        state_byte_0[4]), .C(\state_byte[2]_net_1 ), .Y(
        \state_byte_ns_i_0_0_0[0] ));
    OR3 \state_reset_RNO_1[1]  (.A(\state_reset_ns_i_a2_i_0_0[1] ), .B(
        N_135), .C(\state_reset_RNO_4[1]_net_1 ), .Y(
        \state_reset_ns_i_a2_i_0_2[1] ));
    NOR2A \state_reset_i_RNO_0[0]  (.A(N_174), .B(N_110), .Y(N_150));
    OR2A \state_byte_RNI28611[1]  (.A(size_in[0]), .B(
        \state_byte[1]_net_1 ), .Y(N_64));
    OR3 \state_reset_i_RNO_2[0]  (.A(N_148), .B(N_151), .C(
        \state_reset_ns_i_a2_i_0_0[0] ), .Y(
        \state_reset_ns_i_a2_i_0_2[0] ));
    NOR2 \state_byte_RNITK5G[2]  (.A(\state_byte[2]_net_1 ), .B(
        \state_byte[3]_net_1 ), .Y(N_128));
    DFN1 \state_byte[4]  (.D(\state_byte_nss[4] ), .CLK(FAB_CLK), .Q(
        state_byte_3));
    NOR2A \state_byte_i_RNIKRJ9[0]  (.A(bypass_byte0), .B(
        state_byte_i[0]), .Y(N_118_1));
    MX2 \state_reset_RNO_0[3]  (.A(\state_reset_ns_i_a2_i_0_a7_0_0[3] )
        , .B(N_431), .S(N_110), .Y(N_4));
    NOR2A \state_byte_RNI6C611[3]  (.A(size_in[1]), .B(
        \state_byte[3]_net_1 ), .Y(N_157));
    OR3A \state_byte_i_RNO[0]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        \state_byte_ns[1] ), .C(\state_byte_ns_i_0_0_2[0] ), .Y(
        \state_byte_nss[0] ));
    NOR3B \state_reset_RNO[2]  (.A(N_110), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .C(N_129), .Y(
        \state_reset_nss[2] ));
    AO1 \state_reset_RNO_2[1]  (.A(N_165), .B(N_1006_tz), .C(
        \state_reset_RNO_6[1]_net_1 ), .Y(
        \state_reset_ns_i_a2_i_0_0[1] ));
    DFN1 \state_byte[3]  (.D(\state_byte_nss[3] ), .CLK(FAB_CLK), .Q(
        \state_byte[3]_net_1 ));
    NOR3B \state_reset_i_RNO_9[0]  (.A(size_in[1]), .B(
        \state_byte[3]_net_1 ), .C(size_in[0]), .Y(N_155));
    NOR3C \state_reset_i_RNO_3[0]  (.A(
        \state_reset_ns_i_a2_i_0_a7_0[0] ), .B(N_294), .C(N_95), .Y(
        N_148));
    NOR2B \state_reset_ns_i_a2_i_0_a2_3[1]  (.A(size_in[1]), .B(
        size_in[0]), .Y(N_173));
    NOR2A \state_reset_RNO_0[2]  (.A(N_102), .B(\state_reset[2]_net_1 )
        , .Y(N_129));
    AO1B \state_reset_RNO_9[1]  (.A(\state_reset[3]_net_1 ), .B(
        reset_chain), .C(N_102), .Y(N_1004_tz));
    OR3 \state_reset_RNO_8[1]  (.A(N_430), .B(N_167), .C(
        \state_byte[2]_net_1 ), .Y(N_111));
    VCC VCC_i (.Y(VCC));
    AO1A \state_reset_i_RNO_1[0]  (.A(N_110), .B(
        \state_reset[1]_net_1 ), .C(\state_reset_ns_i_a2_i_0_2[0] ), 
        .Y(\state_reset_ns_i_a2_i_0_3[0] ));
    NOR2A \state_byte_RNISJ5G[1]  (.A(\state_byte[1]_net_1 ), .B(
        \state_byte[3]_net_1 ), .Y(N_176));
    OA1B \state_byte_i_RNIGTTM1[0]  (.A(size_in[0]), .B(size_in[1]), 
        .C(state_byte_i[0]), .Y(\state_byte_ns[1] ));
    DFN1 \state_byte_i[0]  (.D(\state_byte_nss[0] ), .CLK(FAB_CLK), .Q(
        state_byte_i[0]));
    NOR2B \state_byte_RNO[1]  (.A(\state_byte_ns[1] ), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\state_byte_nss[1] ));
    NOR2A \state_byte_RNIV89K2[3]  (.A(\state_byte[3]_net_1 ), .B(N_55)
        , .Y(N_134));
    NOR3B \state_reset_RNO[4]  (.A(N_110), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .C(
        \state_reset_ns_i_a2_0_0_0[4] ), .Y(\state_reset_nss[4] ));
    DFN1 \state_full[1]  (.D(\state_full_nss[1] ), .CLK(FAB_CLK), .Q(
        \state_full[1]_net_1 ));
    OA1B \state_byte_RNI8KC22[3]  (.A(\state_byte[3]_net_1 ), .B(N_166)
        , .C(size_in[1]), .Y(N_167));
    AOI1 \state_reset_RNO_0[4]  (.A(reset_chain), .B(
        \state_reset[3]_net_1 ), .C(\state_reset[4]_net_1 ), .Y(
        \state_reset_ns_i_a2_0_0_0[4] ));
    DFN1 \state_reset_i[0]  (.D(\state_reset_nss[0] ), .CLK(FAB_CLK), 
        .Q(reset_pending));
    OR2 \state_byte_RNIUL5G[2]  (.A(\state_byte[2]_net_1 ), .B(
        state_byte_3), .Y(N_434));
    OR2 \state_reset_RNIS2SS[2]  (.A(\state_reset[2]_net_1 ), .B(
        \state_reset[4]_net_1 ), .Y(N_70));
    NOR3A \state_byte_i_RNIGTTM1_0[0]  (.A(state_byte_i[0]), .B(
        size_in[0]), .C(size_in[1]), .Y(N_159));
    OA1A \state_reset_i_RNINI644[0]  (.A(reset_chain), .B(N_177), .C(
        clear_crc_init_sel_i_0_a7_0), .Y(N_124));
    OA1 \state_reset_RNO[1]  (.A(N_137), .B(
        \state_reset_ns_i_a2_i_0_2[1] ), .C(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\state_reset_nss[1] ));
    DFN1 \state_full[0]  (.D(\state_full_nss[0] ), .CLK(FAB_CLK), .Q(
        \state_full[0]_net_1 ));
    DFN1 \state_reset[3]  (.D(\state_reset_nss[3] ), .CLK(FAB_CLK), .Q(
        \state_reset[3]_net_1 ));
    AO1A \state_full_RNIKV0S5[1]  (.A(N_54), .B(\state_full[1]_net_1 ), 
        .C(N_118), .Y(byte_en));
    XA1 \state_byte_i_RNI0SQR1[0]  (.A(size_in[0]), .B(size_in[1]), .C(
        N_118_1), .Y(N_118));
    NOR3 \state_reset_i_RNO_10[0]  (.A(\state_full[1]_net_1 ), .B(
        reset_pending), .C(N_434), .Y(
        \state_reset_ns_i_a2_i_0_a7_2_0[0] ));
    NOR2B \state_full_RNIK3604[1]  (.A(N_54), .B(\state_full[1]_net_1 )
        , .Y(buffer_full));
    NOR2B \state_byte_RNO[2]  (.A(\state_byte_ns[2] ), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\state_byte_nss[2] ));
    NOR3B \state_full_ns_i_i_0_a7_0[0]  (.A(\state_full[0]_net_1 ), .B(
        N_54), .C(buffer_write_en), .Y(N_146));
    NOR2A \state_byte_RNI28611_0[1]  (.A(\state_byte[1]_net_1 ), .B(
        size_in[0]), .Y(N_166));
    NOR2A \state_reset_RNO_4[1]  (.A(N_1004_tz), .B(N_110), .Y(
        \state_reset_RNO_4[1]_net_1 ));
    OR2A \state_reset_i_RNIA5LN2_0[0]  (.A(reset_chain), .B(
        \state_reset_ns_i_a2_0_0_o2_0[2] ), .Y(N_102));
    AO1 \state_reset_RNO_2[3]  (.A(\state_reset[1]_net_1 ), .B(
        buffer_write_en), .C(N_174), .Y(N_431));
    AO1A \state_full_RNIKV0S5_0[1]  (.A(N_54), .B(
        \state_full[1]_net_1 ), .C(N_118), .Y(byte_en_0));
    DFN1 \state_byte_0[4]  (.D(\state_byte_nss[4] ), .CLK(FAB_CLK), .Q(
        state_byte_0[4]));
    NOR3B \state_reset_i_RNO_8[0]  (.A(size_in[0]), .B(N_176), .C(
        size_in[1]), .Y(N_154));
    OA1 \state_reset_i_RNO_4[0]  (.A(N_154), .B(N_155), .C(
        \state_reset_ns_i_a2_i_0_a7_2_0[0] ), .Y(N_151));
    AO1 \state_reset_RNO_11[1]  (.A(N_438), .B(size_in[1]), .C(
        \state_reset_ns_i_a2_i_0_a7_7_0[1] ), .Y(
        state_reset_ns_i_a2_i_0_125_tz_0));
    NOR2A \state_reset_RNIGROJ2[1]  (.A(\state_reset[1]_net_1 ), .B(
        buffer_write_en), .Y(N_169));
    NOR3A \state_reset_i_RNO_11[0]  (.A(
        \state_reset_ns_i_a2_i_0_a7_4_0[0] ), .B(size_in[0]), .C(
        size_in[1]), .Y(N_153));
    OR2A \state_byte_RNI8KC22[1]  (.A(N_64), .B(N_157), .Y(N_430));
    OR3A \state_byte_0_RNIJLMD9[4]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), 
        .B(N_133), .C(\state_byte_ns_0_0_0_0[4] ), .Y(
        \state_byte_nss[4] ));
    GND GND_i (.Y(GND));
    OR2B state_full_s3_i_i_o2_i_o2 (.A(\state_full[0]_net_1 ), .B(
        \state_full[1]_net_1 ), .Y(bypass_byte0));
    NOR2B \state_byte_RNO[3]  (.A(\state_byte[2]_net_1 ), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\state_byte_nss[3] ));
    OR2 \state_byte_i_RNIOHAP3[0]  (.A(N_159), .B(N_430), .Y(N_54));
    OA1 \state_full_ns_0_i_i_a7[1]  (.A(buffer_write_en), .B(N_54), .C(
        \state_full[1]_net_1 ), .Y(N_122));
    OA1A \state_byte_RNI9P9Q1[1]  (.A(size_in[0]), .B(size_in[1]), .C(
        \state_byte[1]_net_1 ), .Y(\state_byte_ns[2] ));
    DFN1 \state_reset[4]  (.D(\state_reset_nss[4] ), .CLK(FAB_CLK), .Q(
        \state_reset[4]_net_1 ));
    AO1A \state_full_ns_i_i_0_1[0]  (.A(N_54), .B(N_55), .C(
        \state_full_ns_i_i_0_0[0]_net_1 ), .Y(
        \state_full_ns_i_i_0_1[0]_net_1 ));
    NOR3A \state_reset_i_RNO[0]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_150), .C(\state_reset_ns_i_a2_i_0_3[0] ), .Y(
        \state_reset_nss[0] ));
    NOR3 \state_reset_RNI93AB1[4]  (.A(\state_reset[4]_net_1 ), .B(
        \state_reset[3]_net_1 ), .C(\state_reset[1]_net_1 ), .Y(
        clear_crc_init_sel_i_0_a7_0));
    AOI1B \state_byte_RNIJV8A6[4]  (.A(reset_chain), .B(state_byte_3), 
        .C(N_54), .Y(N_125));
    NOR3A \state_reset_i_RNIA5LN2[0]  (.A(reset_chain), .B(
        \state_full[1]_net_1 ), .C(reset_pending), .Y(N_165));
    OA1 \state_reset_RNO_6[1]  (.A(N_173), .B(state_byte_0[4]), .C(
        N_169), .Y(\state_reset_RNO_6[1]_net_1 ));
    NOR3C \state_reset_RNO_10[1]  (.A(size_in[0]), .B(
        \state_byte[1]_net_1 ), .C(state_byte_3), .Y(
        \state_reset_ns_i_a2_i_0_a7_8_0[1] ));
    NOR3A \state_byte_i_RNID47B4[0]  (.A(N_435), .B(size_in[1]), .C(
        N_55), .Y(N_133));
    NOR2B \state_reset_RNO[3]  (.A(N_4), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\state_reset_nss[3] ));
    OA1 \state_reset_RNO_3[1]  (.A(N_169), .B(N_160), .C(N_111), .Y(
        N_135));
    OR3 \state_byte_RNIQU576[3]  (.A(N_430), .B(N_167), .C(
        \state_reset_ns_i_a2_i_0_o2_1_0[3] ), .Y(N_110));
    NOR2A \state_full_RNIOVG56[1]  (.A(buffer_write_en), .B(
        buffer_full), .Y(buffer_en));
    OR2 \state_byte_RNIAMC22[2]  (.A(N_434), .B(N_173), .Y(
        \state_reset_ns_i_a2_i_0_o2_1_0[3] ));
    DFN1 \state_byte[2]  (.D(\state_byte_nss[2] ), .CLK(FAB_CLK), .Q(
        \state_byte[2]_net_1 ));
    NOR2 \state_byte_RNISJ5G_0[1]  (.A(\state_byte[1]_net_1 ), .B(
        \state_byte[3]_net_1 ), .Y(N_294));
    MX2A \state_byte_i_RNI65T51[0]  (.A(state_byte_i[0]), .B(
        \state_byte[1]_net_1 ), .S(size_in[0]), .Y(N_435));
    OA1 \state_reset_RNO_12[1]  (.A(size_in[0]), .B(size_in[1]), .C(
        \state_byte[2]_net_1 ), .Y(\state_reset_ns_i_a2_i_0_a7_2_0[1] )
        );
    NOR2A \state_reset_RNI9J9N2[3]  (.A(\state_reset[3]_net_1 ), .B(
        reset_chain), .Y(N_174));
    NOR3 \state_reset_i_RNO_6[0]  (.A(\state_full[1]_net_1 ), .B(
        reset_pending), .C(\state_byte[2]_net_1 ), .Y(
        \state_reset_ns_i_a2_i_0_a7_0[0] ));
    DFN1 \state_byte[1]  (.D(\state_byte_nss[1] ), .CLK(FAB_CLK), .Q(
        \state_byte[1]_net_1 ));
    OR3 \state_reset_RNO_5[1]  (.A(\state_reset_ns_i_a2_i_0_a7_8_0[1] )
        , .B(state_reset_ns_i_a2_i_0_125_tz_0), .C(
        \state_reset_ns_i_a2_i_0_a7_2_0[1] ), .Y(N_1006_tz));
    NOR2A \state_reset_i_RNIJT0G[0]  (.A(reset_pending), .B(
        state_byte_3), .Y(N_177));
    OR3A \state_byte_i_RNO_0[0]  (.A(N_55), .B(
        \state_byte_ns_i_0_0_0[0] ), .C(\state_byte_ns[2] ), .Y(
        \state_byte_ns_i_0_0_2[0] ));
    DFN1 \state_reset[1]  (.D(\state_reset_nss[1] ), .CLK(FAB_CLK), .Q(
        \state_reset[1]_net_1 ));
    NOR3A \state_reset_i_RNO_12[0]  (.A(state_byte_0[4]), .B(
        \state_full[1]_net_1 ), .C(reset_pending), .Y(
        \state_reset_ns_i_a2_i_0_a7_4_0[0] ));
    OA1 \state_full_srsts[0]  (.A(N_146), .B(
        \state_full_ns_i_i_0_1[0]_net_1 ), .C(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\state_full_nss[0] ));
    AO1A \state_byte_0_RNIIPQV4[4]  (.A(buffer_write_en), .B(
        state_byte_0[4]), .C(N_134), .Y(\state_byte_ns_0_0_0_0[4] ));
    AO1D \state_reset_i_RNO_7[0]  (.A(size_in[1]), .B(size_in[0]), .C(
        state_byte_0[4]), .Y(N_95));
    AO1 \state_reset_RNO_13[1]  (.A(\state_byte[3]_net_1 ), .B(
        state_byte_0[4]), .C(N_176), .Y(N_438));
    AO1D \state_reset_i_RNO_5[0]  (.A(reset_pending), .B(reset_chain), 
        .C(N_153), .Y(\state_reset_ns_i_a2_i_0_0[0] ));
    AXOI7 \state_full_ns_i_i_0_0[0]  (.A(buffer_write_en), .B(
        \state_full[1]_net_1 ), .C(\state_full[0]_net_1 ), .Y(
        \state_full_ns_i_i_0_0[0]_net_1 ));
    NOR2A \state_full_RNIOVG56_0[1]  (.A(buffer_write_en), .B(
        buffer_full), .Y(buffer_en_0));
    OR2 \state_full_RNI0E6C2[1]  (.A(\state_full[1]_net_1 ), .B(
        buffer_write_en), .Y(N_55));
    NOR3A \state_reset_RNO_0[1]  (.A(N_70), .B(buffer_write_en), .C(
        N_110), .Y(N_137));
    DFN1 \state_reset[2]  (.D(\state_reset_nss[2] ), .CLK(FAB_CLK), .Q(
        \state_reset[2]_net_1 ));
    OA1 \state_full_srsts[1]  (.A(N_122), .B(N_123), .C(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\state_full_nss[1] ));
    
endmodule


module bit_reversal_32s_0_1_2_3_4s(
       rev_in_type_0,
       rev_in_type,
       bus_wr_0,
       bus_wr_16,
       bus_wr_1,
       bus_wr_25,
       bus_wr_2,
       bus_wr_3,
       bus_reversed,
       N_358,
       N_350,
       N_351,
       N_337,
       N_366,
       N_367,
       N_357,
       N_349,
       N_352,
       N_360,
       N_336,
       N_365,
       N_356,
       N_348,
       N_353,
       N_361,
       N_335,
       N_364,
       N_332,
       N_355,
       N_362,
       N_334,
       N_333,
       N_363,
       N_347,
       N_354
    );
input  [0:0] rev_in_type_0;
input  [1:0] rev_in_type;
input  bus_wr_0;
input  bus_wr_16;
input  bus_wr_1;
input  bus_wr_25;
input  bus_wr_2;
input  bus_wr_3;
output [31:0] bus_reversed;
input  N_358;
input  N_350;
input  N_351;
input  N_337;
input  N_366;
input  N_367;
input  N_357;
input  N_349;
input  N_352;
input  N_360;
input  N_336;
input  N_365;
input  N_356;
input  N_348;
input  N_353;
input  N_361;
input  N_335;
input  N_364;
input  N_332;
input  N_355;
input  N_362;
input  N_334;
input  N_333;
input  N_363;
input  N_347;
input  N_354;

    wire N_9, N_16, N_24, N_25, N_32, N_33, N_40, N_41, N_48, N_56, 
        N_57, N_64, N_65, N_72, N_10, N_15, N_18, N_26, N_34, N_42, 
        N_47, N_50, N_58, N_66, N_11, N_14, N_19, N_22, N_27, N_30, 
        N_35, N_38, N_43, N_46, N_51, N_54, N_59, N_62, N_67, N_70, 
        N_12, N_28, N_36, N_37, N_44, N_68, N_69, N_60, N_17, N_49, 
        N_23, N_55, N_20, N_52, N_13, N_45, N_39, N_71, N_31, N_63, 
        N_21, N_53, N_29, N_61, GND, VCC;
    
    MX2 \data_out_2[6]  (.A(bus_wr_1), .B(bus_wr_25), .S(
        rev_in_type[1]), .Y(N_47));
    MX2 \data_out_1[3]  (.A(bus_wr_3), .B(N_355), .S(rev_in_type[1]), 
        .Y(N_12));
    MX2 \data_out_3[23]  (.A(N_32), .B(N_64), .S(rev_in_type[0]), .Y(
        bus_reversed[23]));
    MX2 \data_out_1[30]  (.A(N_336), .B(N_360), .S(rev_in_type[1]), .Y(
        N_39));
    MX2 \data_out_3[9]  (.A(N_18), .B(N_50), .S(rev_in_type_0[0]), .Y(
        bus_reversed[9]));
    MX2 \data_out_2[18]  (.A(N_364), .B(N_356), .S(rev_in_type[1]), .Y(
        N_59));
    MX2 \data_out_2[24]  (.A(N_337), .B(N_350), .S(rev_in_type[1]), .Y(
        N_65));
    MX2 \data_out_1[4]  (.A(N_347), .B(N_354), .S(rev_in_type[1]), .Y(
        N_13));
    MX2 \data_out_1[14]  (.A(N_357), .B(bus_wr_1), .S(rev_in_type[1]), 
        .Y(N_23));
    MX2 \data_out_3[15]  (.A(N_24), .B(N_56), .S(rev_in_type_0[0]), .Y(
        bus_reversed[15]));
    MX2 \data_out_1[24]  (.A(N_367), .B(N_366), .S(rev_in_type[1]), .Y(
        N_33));
    MX2 \data_out_1[0]  (.A(bus_wr_0), .B(N_358), .S(rev_in_type[1]), 
        .Y(N_9));
    MX2 \data_out_1[6]  (.A(N_349), .B(N_352), .S(rev_in_type[1]), .Y(
        N_15));
    MX2 \data_out_3[24]  (.A(N_33), .B(N_65), .S(rev_in_type[0]), .Y(
        bus_reversed[24]));
    MX2 \data_out_3[0]  (.A(N_9), .B(N_41), .S(rev_in_type_0[0]), .Y(
        bus_reversed[0]));
    MX2 \data_out_2[28]  (.A(N_333), .B(bus_wr_3), .S(rev_in_type[1]), 
        .Y(N_69));
    MX2 \data_out_2[15]  (.A(N_351), .B(bus_wr_16), .S(rev_in_type[1]), 
        .Y(N_56));
    MX2 \data_out_1[18]  (.A(N_361), .B(N_335), .S(rev_in_type[1]), .Y(
        N_27));
    MX2 \data_out_1[28]  (.A(N_334), .B(N_362), .S(rev_in_type[1]), .Y(
        N_37));
    VCC VCC_i (.Y(VCC));
    MX2 \data_out_3[17]  (.A(N_26), .B(N_58), .S(rev_in_type[0]), .Y(
        bus_reversed[17]));
    MX2 \data_out_2[4]  (.A(bus_wr_3), .B(N_333), .S(rev_in_type[1]), 
        .Y(N_45));
    MX2 \data_out_3[28]  (.A(N_37), .B(N_69), .S(rev_in_type[0]), .Y(
        bus_reversed[28]));
    MX2 \data_out_1[8]  (.A(N_351), .B(N_350), .S(rev_in_type[1]), .Y(
        N_17));
    MX2 \data_out_3[1]  (.A(N_10), .B(N_42), .S(rev_in_type_0[0]), .Y(
        bus_reversed[1]));
    MX2 \data_out_2[8]  (.A(N_358), .B(N_366), .S(rev_in_type[1]), .Y(
        N_49));
    MX2 \data_out_3[16]  (.A(N_25), .B(N_57), .S(rev_in_type[0]), .Y(
        bus_reversed[16]));
    MX2 \data_out_2[17]  (.A(N_365), .B(N_357), .S(rev_in_type[1]), .Y(
        N_58));
    MX2 \data_out_2[25]  (.A(N_336), .B(N_349), .S(rev_in_type[1]), .Y(
        N_66));
    MX2 \data_out_1[15]  (.A(N_358), .B(bus_wr_0), .S(rev_in_type[1]), 
        .Y(N_24));
    MX2 \data_out_3[11]  (.A(N_20), .B(N_52), .S(rev_in_type_0[0]), .Y(
        bus_reversed[11]));
    MX2 \data_out_2[3]  (.A(N_347), .B(N_334), .S(rev_in_type[1]), .Y(
        N_44));
    MX2 \data_out_1[25]  (.A(bus_wr_25), .B(N_365), .S(rev_in_type[1]), 
        .Y(N_34));
    MX2 \data_out_2[2]  (.A(N_348), .B(N_335), .S(rev_in_type[1]), .Y(
        N_43));
    MX2 \data_out_3[3]  (.A(N_12), .B(N_44), .S(rev_in_type_0[0]), .Y(
        bus_reversed[3]));
    MX2 \data_out_3[25]  (.A(N_34), .B(N_66), .S(rev_in_type[0]), .Y(
        bus_reversed[25]));
    MX2 \data_out_2[16]  (.A(N_366), .B(N_358), .S(rev_in_type[1]), .Y(
        N_57));
    MX2 \data_out_3[10]  (.A(N_19), .B(N_51), .S(rev_in_type_0[0]), .Y(
        bus_reversed[10]));
    MX2 \data_out_2[11]  (.A(N_355), .B(N_363), .S(rev_in_type[1]), .Y(
        N_52));
    MX2 \data_out_2[5]  (.A(bus_wr_2), .B(N_332), .S(rev_in_type[1]), 
        .Y(N_46));
    MX2 \data_out_2[27]  (.A(N_334), .B(N_347), .S(rev_in_type[1]), .Y(
        N_68));
    MX2 \data_out_1[17]  (.A(N_360), .B(N_336), .S(rev_in_type[1]), .Y(
        N_26));
    MX2 \data_out_3[12]  (.A(N_21), .B(N_53), .S(rev_in_type_0[0]), .Y(
        bus_reversed[12]));
    MX2 \data_out_1[27]  (.A(N_333), .B(N_363), .S(rev_in_type[1]), .Y(
        N_36));
    MX2 \data_out_2[10]  (.A(N_356), .B(N_364), .S(rev_in_type[1]), .Y(
        N_51));
    MX2 \data_out_3[27]  (.A(N_36), .B(N_68), .S(rev_in_type[0]), .Y(
        bus_reversed[27]));
    MX2 \data_out_2[26]  (.A(N_335), .B(N_348), .S(rev_in_type[1]), .Y(
        N_67));
    MX2 \data_out_1[16]  (.A(bus_wr_16), .B(N_337), .S(rev_in_type[1]), 
        .Y(N_25));
    MX2 \data_out_3[4]  (.A(N_13), .B(N_45), .S(rev_in_type_0[0]), .Y(
        bus_reversed[4]));
    MX2 \data_out_2[12]  (.A(N_354), .B(N_362), .S(rev_in_type[1]), .Y(
        N_53));
    MX2 \data_out_1[26]  (.A(N_332), .B(N_364), .S(rev_in_type[1]), .Y(
        N_35));
    MX2 \data_out_1[1]  (.A(bus_wr_1), .B(N_357), .S(rev_in_type[1]), 
        .Y(N_10));
    GND GND_i (.Y(GND));
    MX2 \data_out_2[21]  (.A(N_361), .B(N_353), .S(rev_in_type[1]), .Y(
        N_62));
    MX2 \data_out_1[7]  (.A(N_350), .B(N_351), .S(rev_in_type[1]), .Y(
        N_16));
    MX2 \data_out_1[11]  (.A(N_354), .B(N_347), .S(rev_in_type[1]), .Y(
        N_20));
    MX2 \data_out_1[9]  (.A(N_352), .B(N_349), .S(rev_in_type[1]), .Y(
        N_18));
    MX2 \data_out_1[21]  (.A(N_364), .B(N_332), .S(rev_in_type[1]), .Y(
        N_30));
    MX2 \data_out_3[26]  (.A(N_35), .B(N_67), .S(rev_in_type[0]), .Y(
        bus_reversed[26]));
    MX2 \data_out_3[21]  (.A(N_30), .B(N_62), .S(rev_in_type[0]), .Y(
        bus_reversed[21]));
    MX2 \data_out_3[19]  (.A(N_28), .B(N_60), .S(rev_in_type[0]), .Y(
        bus_reversed[19]));
    MX2 \data_out_2[20]  (.A(N_362), .B(N_354), .S(rev_in_type[1]), .Y(
        N_61));
    MX2 \data_out_1[10]  (.A(N_353), .B(N_348), .S(rev_in_type[1]), .Y(
        N_19));
    MX2 \data_out_2[9]  (.A(N_357), .B(N_365), .S(rev_in_type[1]), .Y(
        N_50));
    MX2 \data_out_1[20]  (.A(N_363), .B(N_333), .S(rev_in_type[1]), .Y(
        N_29));
    MX2 \data_out_2[7]  (.A(bus_wr_0), .B(N_367), .S(rev_in_type[1]), 
        .Y(N_48));
    MX2 \data_out_2[1]  (.A(N_349), .B(N_336), .S(rev_in_type[1]), .Y(
        N_42));
    MX2 \data_out_2[22]  (.A(N_360), .B(N_352), .S(rev_in_type[1]), .Y(
        N_63));
    MX2 \data_out_1[12]  (.A(N_355), .B(bus_wr_3), .S(rev_in_type[1]), 
        .Y(N_21));
    MX2 \data_out_3[20]  (.A(N_29), .B(N_61), .S(rev_in_type[0]), .Y(
        bus_reversed[20]));
    MX2 \data_out_1[5]  (.A(N_348), .B(N_353), .S(rev_in_type[1]), .Y(
        N_14));
    MX2 \data_out_1[22]  (.A(N_365), .B(bus_wr_25), .S(rev_in_type[1]), 
        .Y(N_31));
    MX2 \data_out_2[19]  (.A(N_363), .B(N_355), .S(rev_in_type[1]), .Y(
        N_60));
    MX2 \data_out_3[8]  (.A(N_17), .B(N_49), .S(rev_in_type_0[0]), .Y(
        bus_reversed[8]));
    MX2 \data_out_2[31]  (.A(N_367), .B(bus_wr_0), .S(rev_in_type[1]), 
        .Y(N_72));
    MX2 \data_out_3[22]  (.A(N_31), .B(N_63), .S(rev_in_type[0]), .Y(
        bus_reversed[22]));
    MX2 \data_out_3[5]  (.A(N_14), .B(N_46), .S(rev_in_type_0[0]), .Y(
        bus_reversed[5]));
    MX2 \data_out_1[2]  (.A(bus_wr_2), .B(N_356), .S(rev_in_type[1]), 
        .Y(N_11));
    MX2 \data_out_3[13]  (.A(N_22), .B(N_54), .S(rev_in_type_0[0]), .Y(
        bus_reversed[13]));
    MX2 \data_out_2[30]  (.A(bus_wr_25), .B(bus_wr_1), .S(
        rev_in_type[1]), .Y(N_71));
    MX2 \data_out_2[29]  (.A(N_332), .B(bus_wr_2), .S(rev_in_type[1]), 
        .Y(N_70));
    MX2 \data_out_1[19]  (.A(N_362), .B(N_334), .S(rev_in_type[1]), .Y(
        N_28));
    MX2 \data_out_1[29]  (.A(N_335), .B(N_361), .S(rev_in_type[1]), .Y(
        N_38));
    MX2 \data_out_2[13]  (.A(N_353), .B(N_361), .S(rev_in_type[1]), .Y(
        N_54));
    MX2 \data_out_2[0]  (.A(N_350), .B(N_337), .S(rev_in_type[1]), .Y(
        N_41));
    MX2 \data_out_3[2]  (.A(N_11), .B(N_43), .S(rev_in_type_0[0]), .Y(
        bus_reversed[2]));
    MX2 \data_out_3[7]  (.A(N_16), .B(N_48), .S(rev_in_type_0[0]), .Y(
        bus_reversed[7]));
    MX2 \data_out_3[31]  (.A(N_40), .B(N_72), .S(rev_in_type[0]), .Y(
        bus_reversed[31]));
    MX2 \data_out_3[29]  (.A(N_38), .B(N_70), .S(rev_in_type[0]), .Y(
        bus_reversed[29]));
    MX2 \data_out_3[6]  (.A(N_15), .B(N_47), .S(rev_in_type_0[0]), .Y(
        bus_reversed[6]));
    MX2 \data_out_3[14]  (.A(N_23), .B(N_55), .S(rev_in_type_0[0]), .Y(
        bus_reversed[14]));
    MX2 \data_out_3[30]  (.A(N_39), .B(N_71), .S(rev_in_type[0]), .Y(
        bus_reversed[30]));
    MX2 \data_out_2[23]  (.A(bus_wr_16), .B(N_351), .S(rev_in_type[1]), 
        .Y(N_64));
    MX2 \data_out_1[13]  (.A(N_356), .B(bus_wr_2), .S(rev_in_type[1]), 
        .Y(N_22));
    MX2 \data_out_2[14]  (.A(N_352), .B(N_360), .S(rev_in_type[1]), .Y(
        N_55));
    MX2 \data_out_1[31]  (.A(N_337), .B(bus_wr_16), .S(rev_in_type[1]), 
        .Y(N_40));
    MX2 \data_out_1[23]  (.A(N_366), .B(N_367), .S(rev_in_type[1]), .Y(
        N_32));
    MX2 \data_out_3[18]  (.A(N_27), .B(N_59), .S(rev_in_type[0]), .Y(
        bus_reversed[18]));
    
endmodule


module \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_0 (
       crc_out_1_0,
       un5_crc_init_justified,
       crc_init_justified_1,
       crc_data_in,
       un90_crc_init_justified,
       crc_in_masked,
       crc_init_justified,
       un79_poly_mux_16,
       un79_poly_mux_0,
       un84_poly_mux_16,
       un84_poly_mux_0,
       un89_poly_mux_16,
       un89_poly_mux_0,
       un94_poly_mux_16,
       un94_poly_mux_0,
       un99_poly_mux_16,
       un99_poly_mux_0,
       \crc_comb_out[2]_23 ,
       \crc_comb_out[2]_15 ,
       \crc_comb_out[2]_0 ,
       poly_mux_17,
       poly_mux_25,
       poly_mux_18,
       poly_mux_6,
       poly_mux_7,
       poly_mux_9,
       poly_mux_4,
       poly_mux_2,
       poly_mux_0,
       un104_poly_mux_16,
       un104_poly_mux_0,
       feedback_29,
       feedback_20,
       feedback_12,
       feedback_22,
       feedback_14,
       feedback_15,
       feedback_16,
       feedback_17,
       feedback_18,
       feedback_9,
       feedback_10,
       feedback_11,
       feedback_5,
       feedback_8,
       feedback_2,
       feedback_1,
       feedback_0_d0,
       feedback_6,
       feedback_4,
       feedback_19,
       feedback_3,
       crc_poly_out_11,
       crc_poly_out_14,
       crc_poly_out_7,
       crc_poly_out_4,
       crc_poly_out_0,
       crc_poly_out_3,
       crc_poly_out_2,
       crc_poly_out_5,
       feedback_0_17,
       feedback_0_10,
       feedback_0_0,
       feedback_0_8,
       un109_poly_mux_16,
       un109_poly_mux_0,
       N_170_0,
       N_170,
       N_170_1,
       crc_poly_size_74_0,
       crc_poly_size_77
    );
output [24:24] crc_out_1_0;
input  [30:30] un5_crc_init_justified;
input  [30:30] crc_init_justified_1;
input  [6:6] crc_data_in;
input  [13:13] un90_crc_init_justified;
output [24:24] crc_in_masked;
input  [23:21] crc_init_justified;
input  un79_poly_mux_16;
input  un79_poly_mux_0;
input  un84_poly_mux_16;
input  un84_poly_mux_0;
input  un89_poly_mux_16;
input  un89_poly_mux_0;
input  un94_poly_mux_16;
input  un94_poly_mux_0;
input  un99_poly_mux_16;
input  un99_poly_mux_0;
output \crc_comb_out[2]_23 ;
output \crc_comb_out[2]_15 ;
output \crc_comb_out[2]_0 ;
input  poly_mux_17;
input  poly_mux_25;
input  poly_mux_18;
input  poly_mux_6;
input  poly_mux_7;
input  poly_mux_9;
input  poly_mux_4;
input  poly_mux_2;
input  poly_mux_0;
input  un104_poly_mux_16;
input  un104_poly_mux_0;
input  feedback_29;
input  feedback_20;
input  feedback_12;
input  feedback_22;
output feedback_14;
output feedback_15;
output feedback_16;
output feedback_17;
output feedback_18;
output feedback_9;
output feedback_10;
output feedback_11;
output feedback_5;
output feedback_8;
output feedback_2;
output feedback_1;
output feedback_0_d0;
output feedback_6;
output feedback_4;
output feedback_19;
output feedback_3;
input  crc_poly_out_11;
input  crc_poly_out_14;
input  crc_poly_out_7;
input  crc_poly_out_4;
input  crc_poly_out_0;
input  crc_poly_out_3;
input  crc_poly_out_2;
input  crc_poly_out_5;
output feedback_0_17;
output feedback_0_10;
output feedback_0_0;
output feedback_0_8;
input  un109_poly_mux_16;
input  un109_poly_mux_0;
output N_170_0;
input  N_170;
output N_170_1;
input  crc_poly_size_74_0;
input  crc_poly_size_77;

    wire un2_feedback_0_net_1, \feedback[23]_net_1 , 
        \feedback[15]_net_1 , GND, VCC;
    
    NOR2B \feedback[15]  (.A(poly_mux_9), .B(N_170_1), .Y(
        \feedback[15]_net_1 ));
    NOR2B \feedback[10]  (.A(poly_mux_4), .B(N_170_1), .Y(feedback_8));
    AX1C \crc_out_1_0[24]  (.A(N_170), .B(poly_mux_17), .C(
        crc_init_justified[22]), .Y(crc_out_1_0[24]));
    OA1 \feedback[17]  (.A(un84_poly_mux_16), .B(un84_poly_mux_0), .C(
        N_170_0), .Y(feedback_15));
    NOR3C \feedback[5]  (.A(crc_poly_size_77), .B(crc_poly_out_5), .C(
        N_170_0), .Y(feedback_3));
    NOR3C \feedback[7]  (.A(crc_poly_size_77), .B(crc_poly_out_7), .C(
        N_170_1), .Y(feedback_5));
    VCC VCC_i (.Y(VCC));
    XOR3 \crc_out_1[15]  (.A(feedback_12), .B(
        un90_crc_init_justified[13]), .C(\feedback[15]_net_1 ), .Y(
        \crc_comb_out[2]_15 ));
    NOR2B \feedback[23]  (.A(poly_mux_17), .B(N_170_1), .Y(
        \feedback[23]_net_1 ));
    NOR2B \feedback[8]  (.A(poly_mux_2), .B(N_170_1), .Y(feedback_6));
    AX1D un2_feedback_0 (.A(un5_crc_init_justified[30]), .B(
        crc_init_justified_1[30]), .C(crc_data_in[6]), .Y(
        un2_feedback_0_net_1));
    NOR3C \feedback[14]  (.A(crc_poly_size_77), .B(crc_poly_out_14), 
        .C(N_170_0), .Y(feedback_0_0));
    NOR2B \feedback[12]  (.A(poly_mux_6), .B(N_170_1), .Y(feedback_10));
    NOR3C \feedback[2]  (.A(crc_poly_size_77), .B(crc_poly_out_2), .C(
        N_170_0), .Y(feedback_0_d0));
    OA1 \feedback[21]  (.A(un104_poly_mux_16), .B(un104_poly_mux_0), 
        .C(N_170_0), .Y(feedback_19));
    OA1 \feedback[19]  (.A(un94_poly_mux_16), .B(un94_poly_mux_0), .C(
        N_170_0), .Y(feedback_17));
    XA1B \crc_in_masked[24]  (.A(feedback_22), .B(
        crc_init_justified[23]), .C(crc_poly_size_74_0), .Y(
        crc_in_masked[24]));
    XOR2 un2_feedback_0_0 (.A(un2_feedback_0_net_1), .B(feedback_29), 
        .Y(N_170_0));
    OA1 \feedback[20]  (.A(un99_poly_mux_16), .B(un99_poly_mux_0), .C(
        N_170_0), .Y(feedback_18));
    XOR2 un2_feedback (.A(un2_feedback_0_net_1), .B(feedback_29), .Y(
        N_170_1));
    NOR2B \feedback[6]  (.A(poly_mux_0), .B(N_170_1), .Y(feedback_4));
    GND GND_i (.Y(GND));
    NOR2B \feedback[31]  (.A(poly_mux_25), .B(N_170_1), .Y(
        feedback_0_17));
    NOR2B \feedback[24]  (.A(poly_mux_18), .B(N_170_1), .Y(
        feedback_0_10));
    OA1 \feedback[22]  (.A(un109_poly_mux_16), .B(un109_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_8));
    XOR3 \crc_out_1[23]  (.A(feedback_20), .B(crc_init_justified[21]), 
        .C(\feedback[23]_net_1 ), .Y(\crc_comb_out[2]_23 ));
    NOR2B \feedback[0]  (.A(crc_poly_out_0), .B(N_170_1), .Y(
        \crc_comb_out[2]_0 ));
    NOR3C \feedback[4]  (.A(crc_poly_size_77), .B(crc_poly_out_4), .C(
        N_170_0), .Y(feedback_2));
    NOR2B \feedback[13]  (.A(poly_mux_7), .B(N_170_1), .Y(feedback_11));
    NOR3C \feedback[3]  (.A(crc_poly_size_77), .B(crc_poly_out_3), .C(
        N_170_0), .Y(feedback_1));
    OA1 \feedback[18]  (.A(un89_poly_mux_16), .B(un89_poly_mux_0), .C(
        N_170_0), .Y(feedback_16));
    OA1 \feedback[16]  (.A(un79_poly_mux_16), .B(un79_poly_mux_0), .C(
        N_170_0), .Y(feedback_14));
    NOR3C \feedback[11]  (.A(crc_poly_size_77), .B(crc_poly_out_11), 
        .C(N_170_0), .Y(feedback_9));
    
endmodule


module \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_4 (
       un70_crc_init_justified_16,
       un70_crc_init_justified_0,
       crc_out_1_4_8,
       crc_out_1_4_0,
       un110_crc_init_justified,
       un25_crc_init_justified,
       crc_init_justified_1,
       crc_data_in,
       crc_out_1_3,
       crc_in_masked_0,
       crc_in_masked_9,
       crc_in_masked_8,
       un104_poly_mux_16,
       un104_poly_mux_0,
       \crc_comb_out[6]_0 ,
       \crc_comb_out[6]_24 ,
       \crc_comb_out[5] ,
       un79_poly_mux_16,
       un79_poly_mux_0,
       un89_poly_mux_16,
       un89_poly_mux_0,
       un94_poly_mux_16,
       un94_poly_mux_0,
       un99_poly_mux_16,
       un99_poly_mux_0,
       un109_poly_mux_16,
       un109_poly_mux_0,
       feedback_0_20,
       feedback_0_10,
       feedback_0_7,
       feedback_0_8,
       feedback_0_9,
       feedback_0_3,
       feedback_0_0,
       feedback_0_11,
       feedback_0_1,
       feedback_0_4,
       feedback_0_2,
       un84_poly_mux_16,
       un84_poly_mux_0,
       poly_mux_4,
       poly_mux_24,
       poly_mux_23,
       poly_mux_22,
       poly_mux_21,
       poly_mux_25,
       poly_mux_17,
       poly_mux_18,
       poly_mux_19,
       poly_mux_2,
       poly_mux_0,
       poly_mux_9,
       poly_mux_7,
       poly_mux_3,
       feedback_29,
       feedback_19,
       feedback_20,
       feedback_17,
       feedback_18,
       feedback_16,
       feedback_11,
       feedback_12,
       feedback_9,
       feedback_10,
       feedback_13,
       feedback_22,
       feedback_25,
       feedback_27,
       feedback_21,
       feedback_23,
       feedback_14,
       feedback_5,
       feedback_6,
       feedback_3,
       feedback_1,
       feedback_2,
       feedback_4,
       feedback_8,
       feedback_15,
       feedback_7,
       feedback_0_d0,
       crc_poly_out_0,
       crc_poly_out_14,
       crc_poly_out_7,
       crc_poly_out_5,
       crc_poly_out_11,
       crc_poly_out_3,
       crc_poly_out_4,
       crc_poly_out_12,
       crc_poly_out_10,
       crc_poly_out_2,
       N_170_0,
       N_170_0_0,
       N_170_0_1,
       N_170,
       N_170_0_2,
       N_170_1,
       crc_poly_size_76_1,
       crc_poly_size_74_0,
       crc_poly_size_75_0,
       crc_poly_size_77
    );
input  un70_crc_init_justified_16;
input  un70_crc_init_justified_0;
output crc_out_1_4_8;
output crc_out_1_4_0;
input  [9:9] un110_crc_init_justified;
input  [26:26] un25_crc_init_justified;
input  [26:26] crc_init_justified_1;
input  [2:2] crc_data_in;
input  [15:15] crc_out_1_3;
output crc_in_masked_0;
output crc_in_masked_9;
input  crc_in_masked_8;
input  un104_poly_mux_16;
input  un104_poly_mux_0;
output \crc_comb_out[6]_0 ;
output \crc_comb_out[6]_24 ;
input  [23:23] \crc_comb_out[5] ;
input  un79_poly_mux_16;
input  un79_poly_mux_0;
input  un89_poly_mux_16;
input  un89_poly_mux_0;
input  un94_poly_mux_16;
input  un94_poly_mux_0;
input  un99_poly_mux_16;
input  un99_poly_mux_0;
input  un109_poly_mux_16;
input  un109_poly_mux_0;
output feedback_0_20;
output feedback_0_10;
output feedback_0_7;
output feedback_0_8;
output feedback_0_9;
output feedback_0_3;
output feedback_0_0;
output feedback_0_11;
output feedback_0_1;
output feedback_0_4;
output feedback_0_2;
input  un84_poly_mux_16;
input  un84_poly_mux_0;
input  poly_mux_4;
input  poly_mux_24;
input  poly_mux_23;
input  poly_mux_22;
input  poly_mux_21;
input  poly_mux_25;
input  poly_mux_17;
input  poly_mux_18;
input  poly_mux_19;
input  poly_mux_2;
input  poly_mux_0;
input  poly_mux_9;
input  poly_mux_7;
input  poly_mux_3;
input  feedback_29;
input  feedback_19;
input  feedback_20;
input  feedback_17;
input  feedback_18;
input  feedback_16;
input  feedback_11;
input  feedback_12;
input  feedback_9;
input  feedback_10;
input  feedback_13;
input  feedback_22;
output feedback_25;
output feedback_27;
output feedback_21;
output feedback_23;
output feedback_14;
output feedback_5;
output feedback_6;
output feedback_3;
output feedback_1;
output feedback_2;
output feedback_4;
output feedback_8;
output feedback_15;
output feedback_7;
output feedback_0_d0;
input  crc_poly_out_0;
input  crc_poly_out_14;
input  crc_poly_out_7;
input  crc_poly_out_5;
input  crc_poly_out_11;
input  crc_poly_out_3;
input  crc_poly_out_4;
input  crc_poly_out_12;
input  crc_poly_out_10;
input  crc_poly_out_2;
output N_170_0;
input  N_170_0_0;
input  N_170_0_1;
input  N_170;
input  N_170_0_2;
output N_170_1;
input  crc_poly_size_76_1;
input  crc_poly_size_74_0;
input  crc_poly_size_75_0;
input  crc_poly_size_77;

    wire un2_feedback_4_net_1, \crc_out_1_2[23]_net_1 , 
        \crc_out_1_0[23]_net_1 , \crc_out_1_2[15]_net_1 , 
        \crc_out_1_0[15]_net_1 , un2_feedback_3_net_1, 
        un2_feedback_2_net_1, un2_feedback_1_net_1, 
        un2_feedback_0_net_1, \feedback_0[24] , GND, VCC;
    
    NOR2B \feedback[15]  (.A(poly_mux_9), .B(N_170_1), .Y(feedback_0_4)
        );
    XOR3 \crc_out_1_2[23]  (.A(feedback_17), .B(
        \crc_out_1_0[23]_net_1 ), .C(feedback_18), .Y(
        \crc_out_1_2[23]_net_1 ));
    NOR2B \feedback[10]  (.A(crc_poly_out_10), .B(N_170_1), .Y(
        feedback_8));
    XOR3 \crc_out_1_4[23]  (.A(feedback_19), .B(
        \crc_out_1_2[23]_net_1 ), .C(feedback_20), .Y(crc_out_1_4_8));
    OA1 \feedback[17]  (.A(un84_poly_mux_16), .B(un84_poly_mux_0), .C(
        N_170_0), .Y(feedback_15));
    NOR3C \feedback[5]  (.A(crc_poly_size_77), .B(crc_poly_out_5), .C(
        N_170_0), .Y(feedback_3));
    AX1D \crc_out_1_0[23]  (.A(un70_crc_init_justified_16), .B(
        un70_crc_init_justified_0), .C(feedback_16), .Y(
        \crc_out_1_0[23]_net_1 ));
    NOR3C \feedback[7]  (.A(crc_poly_size_77), .B(crc_poly_out_7), .C(
        N_170_0), .Y(feedback_5));
    VCC VCC_i (.Y(VCC));
    XOR3 \crc_out_1_2[15]  (.A(feedback_9), .B(\crc_out_1_0[15]_net_1 )
        , .C(feedback_10), .Y(\crc_out_1_2[15]_net_1 ));
    NOR2B \feedback[23]  (.A(poly_mux_17), .B(N_170_1), .Y(feedback_21)
        );
    XOR3 \crc_out_1_4[15]  (.A(feedback_11), .B(
        \crc_out_1_2[15]_net_1 ), .C(feedback_12), .Y(crc_out_1_4_0));
    AX1C un2_feedback_1 (.A(N_170_0_0), .B(poly_mux_21), .C(
        un2_feedback_0_net_1), .Y(un2_feedback_1_net_1));
    NOR2B \feedback[8]  (.A(poly_mux_2), .B(N_170_1), .Y(feedback_6));
    AX1D un2_feedback_0 (.A(un25_crc_init_justified[26]), .B(
        crc_init_justified_1[26]), .C(crc_data_in[2]), .Y(
        un2_feedback_0_net_1));
    NOR3C \feedback[14]  (.A(crc_poly_size_77), .B(crc_poly_out_14), 
        .C(N_170_0), .Y(feedback_0_3));
    AX1C \crc_out_1_0[15]  (.A(N_170_0_0), .B(poly_mux_4), .C(
        un110_crc_init_justified[9]), .Y(\crc_out_1_0[15]_net_1 ));
    NOR2B \feedback[12]  (.A(crc_poly_out_12), .B(N_170_1), .Y(
        feedback_0_1));
    NOR3C \feedback[2]  (.A(crc_poly_size_77), .B(crc_poly_out_2), .C(
        N_170_0), .Y(feedback_0_d0));
    OA1 \feedback[21]  (.A(un104_poly_mux_16), .B(un104_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_10));
    OA1 \feedback[19]  (.A(un94_poly_mux_16), .B(un94_poly_mux_0), .C(
        N_170_0), .Y(feedback_0_8));
    XA1B \crc_in_masked[24]  (.A(feedback_22), .B(crc_in_masked_8), .C(
        crc_poly_size_74_0), .Y(crc_in_masked_9));
    XOR2 un2_feedback_0_0 (.A(un2_feedback_4_net_1), .B(feedback_29), 
        .Y(N_170_0));
    NOR2B \feedback[25]  (.A(poly_mux_19), .B(N_170_1), .Y(feedback_23)
        );
    NOR2B \feedback[9]  (.A(poly_mux_3), .B(N_170_1), .Y(feedback_7));
    AX1C un2_feedback_2 (.A(N_170_0_2), .B(poly_mux_22), .C(
        un2_feedback_1_net_1), .Y(un2_feedback_2_net_1));
    OA1 \feedback[20]  (.A(un99_poly_mux_16), .B(un99_poly_mux_0), .C(
        N_170_0), .Y(feedback_0_9));
    AX1 \crc_out_1[24]  (.A(crc_poly_size_75_0), .B(
        \crc_comb_out[5] [23]), .C(\feedback_0[24] ), .Y(
        \crc_comb_out[6]_24 ));
    XOR2 un2_feedback (.A(un2_feedback_4_net_1), .B(feedback_29), .Y(
        N_170_1));
    NOR2B \feedback[6]  (.A(poly_mux_0), .B(N_170_1), .Y(feedback_4));
    NOR2B \feedback[27]  (.A(poly_mux_21), .B(N_170_1), .Y(feedback_25)
        );
    GND GND_i (.Y(GND));
    AX1C un2_feedback_4 (.A(N_170_0_1), .B(poly_mux_24), .C(
        un2_feedback_3_net_1), .Y(un2_feedback_4_net_1));
    NOR2B \feedback[31]  (.A(poly_mux_25), .B(N_170_1), .Y(
        feedback_0_20));
    AX1C un2_feedback_3 (.A(N_170), .B(poly_mux_23), .C(
        un2_feedback_2_net_1), .Y(un2_feedback_3_net_1));
    NOR2B \feedback[24]  (.A(poly_mux_18), .B(N_170_1), .Y(
        \feedback_0[24] ));
    OA1 \feedback[22]  (.A(un109_poly_mux_16), .B(un109_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_11));
    NOR2B \feedback[29]  (.A(poly_mux_23), .B(N_170_1), .Y(feedback_27)
        );
    NOR2B \feedback[0]  (.A(crc_poly_out_0), .B(N_170_1), .Y(
        \crc_comb_out[6]_0 ));
    XA1B \crc_in_masked[15]  (.A(feedback_13), .B(crc_out_1_3[15]), .C(
        crc_poly_size_76_1), .Y(crc_in_masked_0));
    NOR3C \feedback[4]  (.A(crc_poly_size_77), .B(crc_poly_out_4), .C(
        N_170_0), .Y(feedback_2));
    NOR2B \feedback[13]  (.A(poly_mux_7), .B(N_170_1), .Y(feedback_0_2)
        );
    NOR3C \feedback[3]  (.A(crc_poly_size_77), .B(crc_poly_out_3), .C(
        N_170_0), .Y(feedback_1));
    OA1 \feedback[18]  (.A(un89_poly_mux_16), .B(un89_poly_mux_0), .C(
        N_170_0), .Y(feedback_0_7));
    OA1 \feedback[16]  (.A(un79_poly_mux_16), .B(un79_poly_mux_0), .C(
        N_170_0), .Y(feedback_14));
    NOR2B \feedback[11]  (.A(crc_poly_out_11), .B(N_170_1), .Y(
        feedback_0_0));
    
endmodule


module \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_3 (
       \crc_comb_out[4] ,
       crc_out_1_3,
       un105_crc_init_justified,
       un65_crc_init_justified_16,
       un65_crc_init_justified_0,
       un20_crc_init_justified,
       crc_init_justified_1,
       crc_data_in,
       crc_in_masked,
       crc_out_1_2_0,
       \crc_comb_out[5]_23 ,
       \crc_comb_out[5]_0 ,
       un104_poly_mux_16,
       un104_poly_mux_0,
       un109_poly_mux_16,
       un109_poly_mux_0,
       un84_poly_mux_16,
       un84_poly_mux_0,
       un89_poly_mux_16,
       un89_poly_mux_0,
       un94_poly_mux_16,
       un94_poly_mux_0,
       un99_poly_mux_16,
       un99_poly_mux_0,
       feedback_0_12,
       feedback_0_20,
       feedback_0_10,
       feedback_0_11,
       feedback_0_8,
       feedback_0_9,
       feedback_0_2,
       feedback_0_3,
       feedback_0_0,
       feedback_0_1,
       crc_poly_out_0,
       crc_poly_out_14,
       crc_poly_out_7,
       crc_poly_out_4,
       crc_poly_out_2,
       crc_poly_out_3,
       crc_poly_out_5,
       crc_poly_out_11,
       crc_poly_out_9,
       un79_poly_mux_16,
       un79_poly_mux_0,
       feedback_29,
       feedback_23,
       feedback_11,
       feedback_12,
       feedback_9,
       feedback_10,
       feedback_18,
       feedback_19,
       feedback_17,
       feedback_20,
       feedback_24,
       feedback_26,
       feedback_22,
       feedback_15,
       feedback_16,
       feedback_13,
       feedback_5,
       feedback_2,
       feedback_0_d0,
       feedback_1,
       feedback_4,
       feedback_3,
       feedback_7,
       feedback_14,
       feedback_6,
       poly_mux_19,
       poly_mux_24,
       poly_mux_23,
       poly_mux_22,
       poly_mux_20,
       poly_mux_25,
       poly_mux_17,
       poly_mux_18,
       poly_mux_7,
       poly_mux_9,
       poly_mux_0,
       poly_mux_6,
       poly_mux_2,
       N_170_0,
       crc_poly_size_74,
       N_170,
       N_170_0_0,
       N_170_0_1,
       N_170_0_2,
       crc_poly_size_75_0,
       crc_poly_size_77
    );
input  [24:24] \crc_comb_out[4] ;
output [15:15] crc_out_1_3;
input  [10:10] un105_crc_init_justified;
input  un65_crc_init_justified_16;
input  un65_crc_init_justified_0;
input  [27:27] un20_crc_init_justified;
input  [27:27] crc_init_justified_1;
input  [3:3] crc_data_in;
output [24:23] crc_in_masked;
input  [23:23] crc_out_1_2_0;
output \crc_comb_out[5]_23 ;
output \crc_comb_out[5]_0 ;
input  un104_poly_mux_16;
input  un104_poly_mux_0;
input  un109_poly_mux_16;
input  un109_poly_mux_0;
input  un84_poly_mux_16;
input  un84_poly_mux_0;
input  un89_poly_mux_16;
input  un89_poly_mux_0;
input  un94_poly_mux_16;
input  un94_poly_mux_0;
input  un99_poly_mux_16;
input  un99_poly_mux_0;
input  feedback_0_12;
output feedback_0_20;
output feedback_0_10;
output feedback_0_11;
output feedback_0_8;
output feedback_0_9;
output feedback_0_2;
output feedback_0_3;
output feedback_0_0;
output feedback_0_1;
input  crc_poly_out_0;
input  crc_poly_out_14;
input  crc_poly_out_7;
input  crc_poly_out_4;
input  crc_poly_out_2;
input  crc_poly_out_3;
input  crc_poly_out_5;
input  crc_poly_out_11;
input  crc_poly_out_9;
input  un79_poly_mux_16;
input  un79_poly_mux_0;
input  feedback_29;
output feedback_23;
input  feedback_11;
input  feedback_12;
input  feedback_9;
input  feedback_10;
input  feedback_18;
input  feedback_19;
input  feedback_17;
input  feedback_20;
output feedback_24;
output feedback_26;
output feedback_22;
output feedback_15;
output feedback_16;
output feedback_13;
output feedback_5;
output feedback_2;
output feedback_0_d0;
output feedback_1;
output feedback_4;
output feedback_3;
output feedback_7;
output feedback_14;
output feedback_6;
input  poly_mux_19;
input  poly_mux_24;
input  poly_mux_23;
input  poly_mux_22;
input  poly_mux_20;
input  poly_mux_25;
input  poly_mux_17;
input  poly_mux_18;
input  poly_mux_7;
input  poly_mux_9;
input  poly_mux_0;
input  poly_mux_6;
input  poly_mux_2;
output N_170_0;
input  crc_poly_size_74;
output N_170;
input  N_170_0_0;
input  N_170_0_1;
input  N_170_0_2;
input  crc_poly_size_75_0;
input  crc_poly_size_77;

    wire un2_feedback_3_net_1, \crc_out_1_1[15]_net_1 , 
        \crc_out_1_2[23]_net_1 , \crc_out_1_0[23]_net_1 , 
        un2_feedback_2_net_1, un2_feedback_1_net_1, 
        un2_feedback_0_net_1, \feedback[23]_net_1 , GND, VCC;
    
    NOR2B \feedback[15]  (.A(poly_mux_9), .B(N_170), .Y(feedback_13));
    XOR3 \crc_out_1_2[23]  (.A(feedback_18), .B(
        \crc_out_1_0[23]_net_1 ), .C(feedback_19), .Y(
        \crc_out_1_2[23]_net_1 ));
    OA1 \feedback[17]  (.A(un84_poly_mux_16), .B(un84_poly_mux_0), .C(
        N_170_0), .Y(feedback_15));
    XOR3 \crc_out_1_3[15]  (.A(feedback_11), .B(
        \crc_out_1_1[15]_net_1 ), .C(feedback_12), .Y(crc_out_1_3[15]));
    NOR3C \feedback[5]  (.A(crc_poly_size_77), .B(crc_poly_out_5), .C(
        N_170_0), .Y(feedback_3));
    XA1B \crc_in_masked[23]  (.A(feedback_0_12), .B(crc_out_1_2_0[23]), 
        .C(crc_poly_size_75_0), .Y(crc_in_masked[23]));
    AX1D \crc_out_1_0[23]  (.A(un65_crc_init_justified_16), .B(
        un65_crc_init_justified_0), .C(feedback_17), .Y(
        \crc_out_1_0[23]_net_1 ));
    NOR3C \feedback[7]  (.A(crc_poly_size_77), .B(crc_poly_out_7), .C(
        N_170_0), .Y(feedback_5));
    VCC VCC_i (.Y(VCC));
    NOR2B \feedback[23]  (.A(poly_mux_17), .B(N_170), .Y(
        \feedback[23]_net_1 ));
    AX1C un2_feedback_1 (.A(N_170_0_2), .B(poly_mux_22), .C(
        un2_feedback_0_net_1), .Y(un2_feedback_1_net_1));
    NOR2B \feedback[8]  (.A(poly_mux_2), .B(N_170), .Y(feedback_6));
    AX1D un2_feedback_0 (.A(un20_crc_init_justified[27]), .B(
        crc_init_justified_1[27]), .C(crc_data_in[3]), .Y(
        un2_feedback_0_net_1));
    NOR2B \feedback[28]  (.A(poly_mux_22), .B(N_170), .Y(feedback_26));
    NOR3C \feedback[14]  (.A(crc_poly_size_77), .B(crc_poly_out_14), 
        .C(N_170_0), .Y(feedback_0_3));
    NOR2B \feedback[26]  (.A(poly_mux_20), .B(N_170), .Y(feedback_24));
    NOR2B \feedback[12]  (.A(poly_mux_6), .B(N_170), .Y(feedback_0_1));
    NOR3C \feedback[2]  (.A(crc_poly_size_77), .B(crc_poly_out_2), .C(
        N_170_0), .Y(feedback_0_d0));
    OA1 \feedback[21]  (.A(un104_poly_mux_16), .B(un104_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_10));
    OA1 \feedback[19]  (.A(un94_poly_mux_16), .B(un94_poly_mux_0), .C(
        N_170_0), .Y(feedback_0_8));
    NOR2A \crc_in_masked[24]  (.A(\crc_comb_out[4] [24]), .B(
        crc_poly_size_74), .Y(crc_in_masked[24]));
    XOR2 un2_feedback_0_0 (.A(un2_feedback_3_net_1), .B(feedback_29), 
        .Y(N_170_0));
    AND2 \feedback[25]  (.A(N_170), .B(poly_mux_19), .Y(feedback_23));
    NOR2B \feedback[9]  (.A(crc_poly_out_9), .B(N_170), .Y(feedback_7));
    AX1C un2_feedback_2 (.A(N_170_0_1), .B(poly_mux_23), .C(
        un2_feedback_1_net_1), .Y(un2_feedback_2_net_1));
    OA1 \feedback[20]  (.A(un99_poly_mux_16), .B(un99_poly_mux_0), .C(
        N_170_0), .Y(feedback_0_9));
    XOR2 un2_feedback (.A(un2_feedback_3_net_1), .B(feedback_29), .Y(
        N_170));
    NOR2B \feedback[6]  (.A(poly_mux_0), .B(N_170), .Y(feedback_4));
    GND GND_i (.Y(GND));
    NOR2B \feedback[31]  (.A(poly_mux_25), .B(N_170), .Y(feedback_0_20)
        );
    AX1C un2_feedback_3 (.A(N_170_0_0), .B(poly_mux_24), .C(
        un2_feedback_2_net_1), .Y(un2_feedback_3_net_1));
    NOR2B \feedback[24]  (.A(poly_mux_18), .B(N_170), .Y(feedback_22));
    OA1 \feedback[22]  (.A(un109_poly_mux_16), .B(un109_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_11));
    XOR3 \crc_out_1[23]  (.A(feedback_20), .B(\crc_out_1_2[23]_net_1 ), 
        .C(\feedback[23]_net_1 ), .Y(\crc_comb_out[5]_23 ));
    NOR2B \feedback[0]  (.A(crc_poly_out_0), .B(N_170), .Y(
        \crc_comb_out[5]_0 ));
    NOR3C \feedback[4]  (.A(crc_poly_size_77), .B(crc_poly_out_4), .C(
        N_170_0), .Y(feedback_2));
    NOR2B \feedback[13]  (.A(poly_mux_7), .B(N_170), .Y(feedback_0_2));
    NOR2B \feedback[3]  (.A(crc_poly_out_3), .B(N_170), .Y(feedback_1));
    OA1 \feedback[18]  (.A(un89_poly_mux_16), .B(un89_poly_mux_0), .C(
        N_170_0), .Y(feedback_16));
    OA1 \feedback[16]  (.A(un79_poly_mux_16), .B(un79_poly_mux_0), .C(
        N_170_0), .Y(feedback_14));
    XOR3 \crc_out_1_1[15]  (.A(feedback_9), .B(
        un105_crc_init_justified[10]), .C(feedback_10), .Y(
        \crc_out_1_1[15]_net_1 ));
    NOR3C \feedback[11]  (.A(crc_poly_size_77), .B(crc_poly_out_11), 
        .C(N_170_0), .Y(feedback_0_0));
    
endmodule


module \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_6 (
       un20_crc_out_16,
       un20_crc_out_0,
       \crc_comb_out[3] ,
       un85_crc_init_justified,
       crc_out_1_4_14,
       un80_crc_init_justified,
       crc_out_1_3_14,
       un130_crc_init_justified,
       \crc_comb_out[1] ,
       crc_out_1_6_14,
       crc_out_1_6_2,
       crc_out_1_6_0,
       crc_out_1_6_3,
       crc_out_1_2_0,
       \crc_comb_out[4]_15 ,
       \crc_comb_out[4]_0 ,
       \crc_comb_out[2]_15 ,
       \crc_comb_out[2]_0 ,
       crc_out_1_1_14,
       crc_in_masked_0_9,
       crc_in_masked_0_0,
       \crc_comb_out[5] ,
       crc_init_justified,
       crc_data_in,
       \crc_comb_out[6]_24 ,
       \crc_comb_out[6]_0 ,
       un15_crc_out_0,
       crc_out_1_0_0,
       crc_in_masked_1_9,
       crc_in_masked_1_0,
       crc_in_masked_2_9,
       crc_in_masked_2_0,
       crc_out_1_5_0,
       crc_in_masked_3,
       feedback_30,
       feedback_24,
       feedback_13,
       feedback_12,
       feedback_11,
       feedback_7,
       feedback_27,
       feedback_28,
       feedback_25,
       feedback_26,
       feedback_19,
       feedback_20,
       feedback_17,
       feedback_18,
       feedback_15,
       feedback_16,
       feedback_10,
       feedback_9,
       feedback_6_d0,
       feedback_5_d0,
       feedback_3_d0,
       feedback_4_d0,
       feedback_2_d0,
       feedback_1_d0,
       feedback_21,
       feedback_23,
       crc_in_masked_9,
       crc_in_masked_0_d0,
       crc_in_masked_8,
       feedback_1_24,
       feedback_1_16,
       feedback_1_17,
       feedback_1_15,
       feedback_1_19,
       feedback_1_18,
       feedback_1_7,
       feedback_1_8,
       feedback_1_10,
       feedback_1_11,
       feedback_1_6,
       feedback_1_2,
       feedback_1_3,
       feedback_1_4,
       feedback_1_1,
       feedback_1_9,
       feedback_1_5,
       feedback_1_0,
       feedback_1_20,
       un104_poly_mux_16,
       un104_poly_mux_0,
       un109_poly_mux_16,
       un109_poly_mux_0,
       feedback_6_2,
       feedback_6_13,
       un79_poly_mux_16,
       un79_poly_mux_0,
       feedback_4_5,
       feedback_4_6,
       feedback_4_3,
       feedback_4_1,
       feedback_4_14,
       feedback_4_15,
       feedback_4_4,
       feedback_4_2,
       feedback_4_23,
       feedback_4_16,
       un89_poly_mux_16,
       un89_poly_mux_0,
       feedback_2_23,
       feedback_2_16,
       feedback_2_14,
       feedback_2_15,
       feedback_2_17,
       feedback_2_6,
       feedback_2_5,
       feedback_2_1,
       feedback_2_7,
       feedback_2_3,
       feedback_2_4,
       feedback_2_2,
       feedback_2_0,
       feedback_2_8,
       feedback_2_9,
       feedback_2_18,
       un99_poly_mux_16,
       un99_poly_mux_0,
       un45_crc_out,
       crc_init_mux_6,
       crc_init_mux_2,
       crc_init_mux_4,
       crc_init_mux_0,
       crc_init_mux_3,
       crc_init_mux_1,
       crc_init_mux_7,
       \crc_comb_out[8]_0 ,
       \crc_comb_out[8]_14 ,
       \crc_comb_out[8]_25 ,
       \crc_comb_out[8]_26 ,
       \crc_comb_out[8]_28 ,
       \crc_comb_out[8]_29 ,
       \crc_comb_out[8]_30 ,
       \crc_comb_out[8]_22 ,
       \crc_comb_out[8]_1 ,
       \crc_comb_out[8]_6 ,
       \crc_comb_out[8]_12 ,
       \crc_comb_out[8]_4 ,
       \crc_comb_out[8]_5 ,
       \crc_comb_out[8]_13 ,
       \crc_comb_out[8]_16 ,
       \crc_comb_out[8]_2 ,
       \crc_comb_out[8]_18 ,
       \crc_comb_out[8]_23 ,
       \crc_comb_out[7]_0 ,
       \crc_comb_out[7]_23 ,
       feedback_0_24,
       feedback_0_25,
       feedback_0_18,
       feedback_0_19,
       feedback_0_16,
       feedback_0_17,
       feedback_0_15,
       feedback_0_20,
       feedback_0_11,
       feedback_0_8,
       feedback_0_7,
       feedback_0_6,
       feedback_0_9,
       feedback_0_10,
       feedback_0_2,
       feedback_0_0,
       feedback_0_3,
       feedback_0_4,
       feedback_0_1,
       feedback_0_5,
       feedback_0_27,
       feedback_0_29,
       feedback_0_12,
       feedback_0_14,
       feedback_0_21,
       feedback_0_23,
       un84_poly_mux_16,
       un84_poly_mux_0,
       poly_mux_8,
       poly_mux_26,
       poly_mux_25,
       poly_mux_24,
       poly_mux_28,
       poly_mux_27,
       poly_mux_14,
       poly_mux_7,
       poly_mux_9,
       poly_mux_5,
       poly_mux_0,
       poly_mux_29,
       poly_mux_12,
       poly_mux_30,
       poly_mux_22,
       poly_mux_23,
       poly_mux_11,
       crc_unit_out_0,
       crc_unit_out_1,
       crc_unit_out_6,
       crc_unit_out_25,
       crc_unit_out_9,
       un94_poly_mux_16,
       un94_poly_mux_0,
       feedback_3_16,
       feedback_3_14,
       feedback_3_15,
       feedback_3_5,
       feedback_3_6,
       feedback_3_3,
       feedback_3_1,
       feedback_3_7,
       feedback_3_4,
       feedback_3_0,
       feedback_3_2,
       feedback_3_23,
       feedback_3_8,
       feedback_3_9,
       crc_poly_out_9,
       crc_poly_out_0,
       crc_poly_out_4,
       crc_poly_out_2,
       crc_poly_out_7,
       crc_poly_out_5,
       crc_poly_out_6,
       crc_poly_out_14,
       crc_poly_out_3,
       crc_poly_out_11,
       feedback_5_5,
       feedback_5_1,
       feedback_5_14,
       feedback_5_0,
       feedback_5_6,
       feedback_5_2,
       N_170_0,
       N_170_0_0,
       N_170_1,
       N_170_2,
       crc_poly_size_74_0,
       N_170_0_1,
       N_170_0_2,
       N_170_0_3,
       N_170_3,
       crc_poly_size_76_0,
       crc_poly_size_77,
       N_170_0_4,
       N_170_4,
       N_170_5,
       N_170_6,
       N_170_0_5,
       N_170_0_6,
       crc_poly_size_76_1,
       crc_poly_size_75_0
    );
input  un20_crc_out_16;
input  un20_crc_out_0;
input  [24:24] \crc_comb_out[3] ;
input  [14:14] un85_crc_init_justified;
output crc_out_1_4_14;
input  [15:15] un80_crc_init_justified;
output crc_out_1_3_14;
input  [5:5] un130_crc_init_justified;
input  [0:0] \crc_comb_out[1] ;
output crc_out_1_6_14;
output crc_out_1_6_2;
output crc_out_1_6_0;
output crc_out_1_6_3;
output crc_out_1_2_0;
input  \crc_comb_out[4]_15 ;
input  \crc_comb_out[4]_0 ;
input  \crc_comb_out[2]_15 ;
input  \crc_comb_out[2]_0 ;
output crc_out_1_1_14;
input  crc_in_masked_0_9;
input  crc_in_masked_0_0;
input  [0:0] \crc_comb_out[5] ;
input  [24:24] crc_init_justified;
input  [0:0] crc_data_in;
input  \crc_comb_out[6]_24 ;
input  \crc_comb_out[6]_0 ;
input  un15_crc_out_0;
input  [3:3] crc_out_1_0_0;
input  crc_in_masked_1_9;
input  crc_in_masked_1_0;
input  crc_in_masked_2_9;
output crc_in_masked_2_0;
input  [15:15] crc_out_1_5_0;
output [24:24] crc_in_masked_3;
input  feedback_30;
input  feedback_24;
input  feedback_13;
input  feedback_12;
input  feedback_11;
input  feedback_7;
input  feedback_27;
input  feedback_28;
input  feedback_25;
input  feedback_26;
input  feedback_19;
input  feedback_20;
input  feedback_17;
input  feedback_18;
input  feedback_15;
input  feedback_16;
input  feedback_10;
input  feedback_9;
input  feedback_6_d0;
input  feedback_5_d0;
input  feedback_3_d0;
input  feedback_4_d0;
input  feedback_2_d0;
input  feedback_1_d0;
input  feedback_21;
input  feedback_23;
input  crc_in_masked_9;
input  crc_in_masked_0_d0;
input  crc_in_masked_8;
input  feedback_1_24;
input  feedback_1_16;
input  feedback_1_17;
input  feedback_1_15;
input  feedback_1_19;
input  feedback_1_18;
input  feedback_1_7;
input  feedback_1_8;
input  feedback_1_10;
input  feedback_1_11;
input  feedback_1_6;
input  feedback_1_2;
input  feedback_1_3;
input  feedback_1_4;
input  feedback_1_1;
input  feedback_1_9;
input  feedback_1_5;
input  feedback_1_0;
output feedback_1_20;
input  un104_poly_mux_16;
input  un104_poly_mux_0;
input  un109_poly_mux_16;
input  un109_poly_mux_0;
input  feedback_6_2;
output feedback_6_13;
input  un79_poly_mux_16;
input  un79_poly_mux_0;
input  feedback_4_5;
input  feedback_4_6;
input  feedback_4_3;
input  feedback_4_1;
input  feedback_4_14;
input  feedback_4_15;
input  feedback_4_4;
input  feedback_4_2;
output feedback_4_23;
output feedback_4_16;
input  un89_poly_mux_16;
input  un89_poly_mux_0;
input  feedback_2_23;
input  feedback_2_16;
input  feedback_2_14;
input  feedback_2_15;
input  feedback_2_17;
input  feedback_2_6;
input  feedback_2_5;
input  feedback_2_1;
input  feedback_2_7;
input  feedback_2_3;
input  feedback_2_4;
input  feedback_2_2;
input  feedback_2_0;
input  feedback_2_8;
input  feedback_2_9;
output feedback_2_18;
input  un99_poly_mux_16;
input  un99_poly_mux_0;
input  [25:25] un45_crc_out;
input  crc_init_mux_6;
input  crc_init_mux_2;
input  crc_init_mux_4;
input  crc_init_mux_0;
input  crc_init_mux_3;
input  crc_init_mux_1;
input  crc_init_mux_7;
output \crc_comb_out[8]_0 ;
output \crc_comb_out[8]_14 ;
output \crc_comb_out[8]_25 ;
output \crc_comb_out[8]_26 ;
output \crc_comb_out[8]_28 ;
output \crc_comb_out[8]_29 ;
output \crc_comb_out[8]_30 ;
output \crc_comb_out[8]_22 ;
output \crc_comb_out[8]_1 ;
output \crc_comb_out[8]_6 ;
output \crc_comb_out[8]_12 ;
output \crc_comb_out[8]_4 ;
output \crc_comb_out[8]_5 ;
output \crc_comb_out[8]_13 ;
output \crc_comb_out[8]_16 ;
output \crc_comb_out[8]_2 ;
output \crc_comb_out[8]_18 ;
output \crc_comb_out[8]_23 ;
input  \crc_comb_out[7]_0 ;
input  \crc_comb_out[7]_23 ;
input  feedback_0_24;
input  feedback_0_25;
input  feedback_0_18;
input  feedback_0_19;
input  feedback_0_16;
input  feedback_0_17;
input  feedback_0_15;
input  feedback_0_20;
input  feedback_0_11;
input  feedback_0_8;
input  feedback_0_7;
input  feedback_0_6;
input  feedback_0_9;
input  feedback_0_10;
input  feedback_0_2;
input  feedback_0_0;
input  feedback_0_3;
input  feedback_0_4;
input  feedback_0_1;
input  feedback_0_5;
input  feedback_0_27;
input  feedback_0_29;
input  feedback_0_12;
input  feedback_0_14;
output feedback_0_21;
output feedback_0_23;
input  un84_poly_mux_16;
input  un84_poly_mux_0;
input  poly_mux_8;
input  poly_mux_26;
input  poly_mux_25;
input  poly_mux_24;
input  poly_mux_28;
input  poly_mux_27;
input  poly_mux_14;
input  poly_mux_7;
input  poly_mux_9;
input  poly_mux_5;
input  poly_mux_0;
input  poly_mux_29;
input  poly_mux_12;
input  poly_mux_30;
input  poly_mux_22;
input  poly_mux_23;
input  poly_mux_11;
output crc_unit_out_0;
output crc_unit_out_1;
output crc_unit_out_6;
output crc_unit_out_25;
output crc_unit_out_9;
input  un94_poly_mux_16;
input  un94_poly_mux_0;
input  feedback_3_16;
input  feedback_3_14;
input  feedback_3_15;
input  feedback_3_5;
input  feedback_3_6;
input  feedback_3_3;
input  feedback_3_1;
input  feedback_3_7;
input  feedback_3_4;
input  feedback_3_0;
input  feedback_3_2;
input  feedback_3_23;
output feedback_3_8;
output feedback_3_9;
input  crc_poly_out_9;
input  crc_poly_out_0;
input  crc_poly_out_4;
input  crc_poly_out_2;
input  crc_poly_out_7;
input  crc_poly_out_5;
input  crc_poly_out_6;
input  crc_poly_out_14;
input  crc_poly_out_3;
input  crc_poly_out_11;
input  feedback_5_5;
input  feedback_5_1;
input  feedback_5_14;
input  feedback_5_0;
output feedback_5_6;
output feedback_5_2;
output N_170_0;
input  N_170_0_0;
input  N_170_1;
input  N_170_2;
input  crc_poly_size_74_0;
input  N_170_0_1;
input  N_170_0_2;
input  N_170_0_3;
input  N_170_3;
input  crc_poly_size_76_0;
input  crc_poly_size_77;
input  N_170_0_4;
input  N_170_4;
input  N_170_5;
input  N_170_6;
input  N_170_0_5;
input  N_170_0_6;
input  crc_poly_size_76_1;
input  crc_poly_size_75_0;

    wire un2_feedback_6_net_1, \feedback[9]_net_1 , N_170, 
        \feedback[1] , \crc_out_1_0[28]_net_1 , 
        \crc_out_1_6[15]_net_1 , \crc_out_1_5[15]_net_1 , 
        \crc_out_1_4[15]_net_1 , \crc_out_1_3[15] , 
        \crc_out_1_6[9]_net_1 , \crc_out_1_5[9] , \feedback[15] , 
        \crc_comb_out[8][9] , \crc_out_1_1[4] , \un20_crc_out[28] , 
        \crc_out_1_4[31]_net_1 , \crc_out_1_2[31]_net_1 , 
        \crc_out_1_1[31]_net_1 , \crc_out_1_0[31]_net_1 , 
        \crc_out_1_2[29]_net_1 , \crc_out_1_0[29]_net_1 , 
        \crc_out_1_4[30]_net_1 , \crc_out_1_3[30]_net_1 , 
        \crc_out_1_2[30]_net_1 , \crc_out_1_1[30]_net_1 , 
        \crc_out_1_0[30]_net_1 , \crc_out_1_2[28] , \crc_out_1_1[28] , 
        \crc_out_1_1[27]_net_1 , \crc_out_1_0[26]_net_1 , 
        \crc_out_1_4[22]_net_1 , \crc_out_1_2[22]_net_1 , 
        \crc_out_1_0[22]_net_1 , \crc_out_1_2[21]_net_1 , 
        \crc_out_1_0[21]_net_1 , \crc_out_1_2[19]_net_1 , 
        \crc_out_1_0[19]_net_1 , \crc_out_1_5[23]_net_1 , 
        \crc_out_1_3[23]_net_1 , \crc_out_1_1[23]_net_1 , 
        \crc_out_1_1[20]_net_1 , \crc_out_1_5[14]_net_1 , 
        \crc_out_1_3[14]_net_1 , \crc_out_1_1[14]_net_1 , 
        \crc_out_1_4[10]_net_1 , \crc_out_1_2[10]_net_1 , 
        \crc_out_1_0[10]_net_1 , \crc_out_1_1[15] , \crc_out_1_0[15] , 
        \un120_crc_init_justified[7] , \crc_out_1_6[13]_net_1 , 
        \crc_out_1_4[13]_net_1 , \crc_out_1_3[13]_net_1 , 
        \crc_out_1_2[13]_net_1 , \crc_out_1_0[13]_net_1 , 
        \crc_out_1_2[5]_net_1 , \crc_out_1_0[5]_net_1 , 
        \crc_out_1_4[7]_net_1 , \crc_out_1_2[7]_net_1 , 
        \crc_out_1_0[7]_net_1 , \crc_out_1_3[9] , \crc_out_1_1[9] , 
        \un150_crc_init_justified[1] , \crc_out_1_5[12]_net_1 , 
        \crc_out_1_3[12]_net_1 , \crc_out_1_1[12]_net_1 , 
        \crc_out_1_4[8]_net_1 , \crc_out_1_2[8]_net_1 , 
        \crc_out_1_0[8]_net_1 , \crc_out_1_4[11]_net_1 , 
        \crc_out_1_2[11]_net_1 , \crc_out_1_0[11]_net_1 , 
        \crc_out_1_0[4]_net_1 , \crc_out_1_3[6]_net_1 , 
        \crc_out_1_1[6]_net_1 , \crc_out_1_0[6]_net_1 , 
        \crc_out_1_0[3]_net_1 , un2_feedback_5_net_1, 
        un2_feedback_4_net_1, un2_feedback_3_net_1, 
        un2_feedback_2_net_1, un2_feedback_1_net_1, \feedback_1[26] , 
        \feedback_0[27] , \feedback_0[29] , \feedback[30]_net_1 , 
        \feedback_0[31] , \feedback[23]_net_1 , \feedback_4[2] , 
        \un15_crc_out[28] , \feedback_6[7] , \feedback_5[5] , 
        \feedback_5[6] , \feedback_0[14] , \feedback_5[17] , 
        \crc_comb_out[8][12] , \feedback_2[12] , \feedback_6[3] , 
        \feedback_3[19] , \feedback_1[28] , \un60_crc_out[28] , GND, 
        VCC;
    
    XOR2 \crc_out_1_6[9]  (.A(feedback_7), .B(\crc_out_1_5[9] ), .Y(
        \crc_out_1_6[9]_net_1 ));
    AX1 \crc_out_1[24]  (.A(crc_poly_size_75_0), .B(
        \crc_comb_out[7]_23 ), .C(feedback_0_23), .Y(
        \crc_comb_out[8]_23 ));
    XOR3 \crc_out_1_4[10]  (.A(feedback_5_d0), .B(
        \crc_out_1_2[10]_net_1 ), .C(feedback_0_6), .Y(
        \crc_out_1_4[10]_net_1 ));
    XOR3 \crc_out_1_2[11]  (.A(feedback_4_3), .B(
        \crc_out_1_0[11]_net_1 ), .C(feedback_3_4), .Y(
        \crc_out_1_2[11]_net_1 ));
    OA1 \feedback[21]  (.A(un104_poly_mux_16), .B(un104_poly_mux_0), 
        .C(N_170_0), .Y(feedback_1_20));
    OA1 \feedback[22]  (.A(un109_poly_mux_16), .B(un109_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_21));
    AX1C \crc_out_1_2[30]  (.A(N_170_0_3), .B(poly_mux_26), .C(
        \crc_out_1_1[30]_net_1 ), .Y(\crc_out_1_2[30]_net_1 ));
    NOR2B \feedback[23]  (.A(poly_mux_22), .B(N_170), .Y(
        \feedback[23]_net_1 ));
    OA1 \feedback[20]  (.A(un99_poly_mux_16), .B(un99_poly_mux_0), .C(
        N_170_0), .Y(feedback_2_18));
    XOR3 \crc_out_1_4[8]  (.A(feedback_2_2), .B(\crc_out_1_2[8]_net_1 )
        , .C(feedback_3_3), .Y(\crc_out_1_4[8]_net_1 ));
    AX1C \crc_out_1_4[13]  (.A(N_170_0_3), .B(poly_mux_9), .C(
        \crc_out_1_3[13]_net_1 ), .Y(\crc_out_1_4[13]_net_1 ));
    XOR2 \crc_out_1[26]  (.A(\crc_out_1_0[26]_net_1 ), .B(
        \feedback_1[26] ), .Y(\crc_comb_out[8]_25 ));
    OA1 \feedback[19]  (.A(un94_poly_mux_16), .B(un94_poly_mux_0), .C(
        N_170_0), .Y(\feedback_3[19] ));
    XOR3 \crc_out_1_2[21]  (.A(feedback_0_16), .B(
        \crc_out_1_0[21]_net_1 ), .C(feedback_0_17), .Y(
        \crc_out_1_2[21]_net_1 ));
    XOR3 \crc_out_1_6[22]  (.A(feedback_19), .B(
        \crc_out_1_4[22]_net_1 ), .C(feedback_20), .Y(crc_out_1_6_14));
    AO1 \crc_out_1_0_RNIVQ47TB2[28]  (.A(\crc_comb_out[8]_28 ), .B(
        crc_poly_size_74_0), .C(\crc_out_1_1[4] ), .Y(crc_unit_out_1));
    XOR2 \crc_out_1[19]  (.A(\crc_out_1_2[19]_net_1 ), .B(
        \feedback_3[19] ), .Y(\crc_comb_out[8]_18 ));
    AX1C \crc_out_1_0[5]  (.A(N_170_1), .B(crc_poly_out_0), .C(
        feedback_0_0), .Y(\crc_out_1_0[5]_net_1 ));
    AX1C un2_feedback_2 (.A(N_170_0_6), .B(poly_mux_25), .C(
        un2_feedback_1_net_1), .Y(un2_feedback_2_net_1));
    NOR2B \feedback[6]  (.A(crc_poly_out_6), .B(N_170), .Y(
        \feedback_5[6] ));
    AX1C \crc_out_1_0[4]  (.A(N_170_4), .B(poly_mux_0), .C(
        \crc_comb_out[4]_0 ), .Y(\crc_out_1_0[4]_net_1 ));
    AO1 \crc_out_1_0_RNIQSUNS21[28]  (.A(\crc_comb_out[8][12] ), .B(
        crc_poly_size_77), .C(\un60_crc_out[28] ), .Y(crc_unit_out_9));
    XOR2 \crc_out_1[30]  (.A(\crc_out_1_4[30]_net_1 ), .B(
        \feedback[30]_net_1 ), .Y(\crc_comb_out[8]_29 ));
    AND2 \feedback[9]  (.A(N_170), .B(poly_mux_8), .Y(
        \feedback[9]_net_1 ));
    AX1C \crc_out_1_3[30]  (.A(N_170_0_2), .B(poly_mux_27), .C(
        \crc_out_1_2[30]_net_1 ), .Y(\crc_out_1_3[30]_net_1 ));
    GND GND_i (.Y(GND));
    OA1 \feedback[16]  (.A(un79_poly_mux_16), .B(un79_poly_mux_0), .C(
        N_170_0), .Y(feedback_6_13));
    XOR3 \crc_out_1_2[8]  (.A(feedback_2_0), .B(\crc_out_1_0[8]_net_1 )
        , .C(feedback_3_1), .Y(\crc_out_1_2[8]_net_1 ));
    NOR2B \crc_out_1_RNO[1]  (.A(poly_mux_0), .B(N_170), .Y(
        \feedback[1] ));
    AO1 \crc_out_1_RNIAH8TRM2[9]  (.A(\crc_comb_out[8][9] ), .B(
        crc_poly_size_77), .C(un45_crc_out[25]), .Y(crc_unit_out_6));
    XA1 \crc_out_1_0_RNIOMSNFC2_1[28]  (.A(\feedback_1[28] ), .B(
        \crc_out_1_2[28] ), .C(crc_poly_size_75_0), .Y(
        \un20_crc_out[28] ));
    AX1C \crc_out_1_0[22]  (.A(N_170_3), .B(poly_mux_14), .C(
        un85_crc_init_justified[14]), .Y(\crc_out_1_0[22]_net_1 ));
    XOR2 \crc_out_1_6[15]  (.A(feedback_13), .B(
        \crc_out_1_5[15]_net_1 ), .Y(\crc_out_1_6[15]_net_1 ));
    XA1 \crc_out_1_0_RNIOMSNFC2_2[28]  (.A(\feedback_1[28] ), .B(
        \crc_out_1_2[28] ), .C(crc_poly_size_76_1), .Y(
        \un60_crc_out[28] ));
    XOR3 \crc_out_1_1[27]  (.A(feedback_1_24), .B(crc_in_masked_2_9), 
        .C(feedback_0_25), .Y(\crc_out_1_1[27]_net_1 ));
    XOR3 \crc_out_1[3]  (.A(feedback_5_0), .B(\crc_out_1_0[3]_net_1 ), 
        .C(\feedback_6[3] ), .Y(\crc_comb_out[8]_2 ));
    XOR3 \crc_out_1_3[14]  (.A(feedback_0_8), .B(
        \crc_out_1_1[14]_net_1 ), .C(feedback_9), .Y(
        \crc_out_1_3[14]_net_1 ));
    XOR3 \crc_out_1[5]  (.A(feedback_4_2), .B(\crc_out_1_2[5]_net_1 ), 
        .C(\feedback_5[5] ), .Y(\crc_comb_out[8]_4 ));
    XOR3 \crc_out_1_3[12]  (.A(feedback_3_5), .B(
        \crc_out_1_1[12]_net_1 ), .C(feedback_3_6), .Y(
        \crc_out_1_3[12]_net_1 ));
    AX1C \crc_out_1_0[10]  (.A(crc_poly_size_77), .B(crc_init_mux_2), 
        .C(feedback_2_d0), .Y(\crc_out_1_0[10]_net_1 ));
    AX1C un2_feedback_3 (.A(N_170_0_5), .B(poly_mux_26), .C(
        un2_feedback_2_net_1), .Y(un2_feedback_3_net_1));
    OA1 \feedback[18]  (.A(un89_poly_mux_16), .B(un89_poly_mux_0), .C(
        N_170_0), .Y(feedback_4_16));
    AX1C \crc_out_1_1[30]  (.A(N_170_0_0), .B(poly_mux_25), .C(
        \crc_out_1_0[30]_net_1 ), .Y(\crc_out_1_1[30]_net_1 ));
    NOR2B \feedback[8]  (.A(poly_mux_7), .B(N_170), .Y(feedback_5_6));
    NOR2B \crc_out_1_4_RNO_2[15]  (.A(crc_init_mux_7), .B(
        crc_poly_size_77), .Y(\un120_crc_init_justified[7] ));
    XOR3 \crc_out_1_2[4]  (.A(feedback_3_0), .B(\crc_out_1_0[4]_net_1 )
        , .C(feedback_4_1), .Y(crc_out_1_2_0));
    VCC VCC_i (.Y(VCC));
    AX1 \crc_out_1_0[26]  (.A(crc_poly_size_74_0), .B(
        \crc_comb_out[6]_24 ), .C(feedback_2_23), .Y(
        \crc_out_1_0[26]_net_1 ));
    XOR2 \crc_out_1[27]  (.A(\crc_out_1_1[27]_net_1 ), .B(
        \feedback_0[27] ), .Y(\crc_comb_out[8]_26 ));
    AX1C \crc_out_1[13]  (.A(N_170_0), .B(poly_mux_12), .C(
        \crc_out_1_6[13]_net_1 ), .Y(\crc_comb_out[8]_12 ));
    XOR3 \crc_out_1_6[10]  (.A(feedback_1_7), .B(
        \crc_out_1_4[10]_net_1 ), .C(feedback_1_8), .Y(crc_out_1_6_2));
    XOR3 \crc_out_1_4[21]  (.A(feedback_0_18), .B(
        \crc_out_1_2[21]_net_1 ), .C(feedback_0_19), .Y(crc_out_1_4_14)
        );
    XOR3 \crc_out_1_4[11]  (.A(feedback_5_5), .B(
        \crc_out_1_2[11]_net_1 ), .C(feedback_4_6), .Y(
        \crc_out_1_4[11]_net_1 ));
    NOR2B \crc_out_1_RNO[15]  (.A(poly_mux_14), .B(N_170), .Y(
        \feedback[15] ));
    NOR2B \feedback[24]  (.A(poly_mux_23), .B(N_170), .Y(feedback_0_23)
        );
    AX1 \crc_out_1_0[19]  (.A(crc_poly_size_76_0), .B(
        \crc_comb_out[4]_15 ), .C(feedback_1_15), .Y(
        \crc_out_1_0[19]_net_1 ));
    XOR3 \crc_out_1[12]  (.A(feedback_2_9), .B(\crc_out_1_5[12]_net_1 )
        , .C(\feedback_2[12] ), .Y(\crc_comb_out[8][12] ));
    XOR3 \crc_out_1_6_RNO[9]  (.A(feedback_0_5), .B(\crc_out_1_3[9] ), 
        .C(feedback_2_5), .Y(\crc_out_1_5[9] ));
    XOR3 \crc_out_1[31]  (.A(feedback_0_29), .B(
        \crc_out_1_4[31]_net_1 ), .C(\feedback_0[31] ), .Y(
        \crc_comb_out[8]_30 ));
    AX1C \crc_out_1_0[13]  (.A(N_170_0_4), .B(poly_mux_5), .C(
        un130_crc_init_justified[5]), .Y(\crc_out_1_0[13]_net_1 ));
    XOR3 \crc_out_1_1[20]  (.A(feedback_3_14), .B(crc_in_masked_0_d0), 
        .C(feedback_3_15), .Y(\crc_out_1_1[20]_net_1 ));
    XOR3 \crc_out_1_4[7]  (.A(feedback_0_3), .B(\crc_out_1_2[7]_net_1 )
        , .C(feedback_0_4), .Y(\crc_out_1_4[7]_net_1 ));
    AX1C \crc_out_1_2[31]  (.A(N_170_0_0), .B(poly_mux_26), .C(
        \crc_out_1_1[31]_net_1 ), .Y(\crc_out_1_2[31]_net_1 ));
    NOR3C \feedback[11]  (.A(crc_poly_size_77), .B(crc_poly_out_11), 
        .C(N_170_0), .Y(feedback_3_9));
    NOR3C \feedback[2]  (.A(crc_poly_size_77), .B(crc_poly_out_2), .C(
        N_170_0), .Y(\feedback_4[2] ));
    NOR2B \feedback[12]  (.A(poly_mux_11), .B(N_170), .Y(
        \feedback_2[12] ));
    NOR2B \feedback[25]  (.A(poly_mux_24), .B(N_170), .Y(feedback_4_23)
        );
    XOR2 \crc_out_1[15]  (.A(\feedback[15] ), .B(
        \crc_out_1_6[15]_net_1 ), .Y(\crc_comb_out[8]_14 ));
    NOR2B \feedback[27]  (.A(poly_mux_26), .B(N_170), .Y(
        \feedback_0[27] ));
    AX1C \crc_out_1_0[30]  (.A(N_170_1), .B(poly_mux_24), .C(
        crc_in_masked_1_9), .Y(\crc_out_1_0[30]_net_1 ));
    XOR3 \crc_out_1[14]  (.A(feedback_0_12), .B(
        \crc_out_1_5[14]_net_1 ), .C(\feedback_0[14] ), .Y(
        \crc_comb_out[8]_13 ));
    NOR2B \feedback[10]  (.A(poly_mux_9), .B(N_170_0), .Y(feedback_3_8)
        );
    XOR3 \crc_out_1_6[13]  (.A(feedback_1_10), .B(
        \crc_out_1_4[13]_net_1 ), .C(feedback_1_11), .Y(
        \crc_out_1_6[13]_net_1 ));
    AX1 \crc_out_1_0[29]  (.A(crc_poly_size_74_0), .B(
        \crc_comb_out[3] [24]), .C(feedback_0_24), .Y(
        \crc_out_1_0[29]_net_1 ));
    XOR3 \crc_out_1[2]  (.A(feedback_1_0), .B(\crc_comb_out[6]_0 ), .C(
        \feedback_4[2] ), .Y(\crc_comb_out[8]_1 ));
    AX1C un2_feedback_5 (.A(N_170_0_3), .B(poly_mux_28), .C(
        un2_feedback_4_net_1), .Y(un2_feedback_5_net_1));
    XOR3 \crc_out_1_1[23]  (.A(feedback_2_14), .B(
        un80_crc_init_justified[15]), .C(feedback_2_15), .Y(
        \crc_out_1_1[23]_net_1 ));
    XOR3 \crc_out_1_3[6]  (.A(feedback_5_1), .B(\crc_out_1_1[6]_net_1 )
        , .C(feedback_3_2), .Y(\crc_out_1_3[6]_net_1 ));
    NOR2B \feedback[31]  (.A(poly_mux_30), .B(N_170), .Y(
        \feedback_0[31] ));
    AX1C \crc_out_1_4[30]  (.A(N_170_0_1), .B(poly_mux_28), .C(
        \crc_out_1_3[30]_net_1 ), .Y(\crc_out_1_4[30]_net_1 ));
    XOR3 \crc_out_1_2[22]  (.A(feedback_15), .B(
        \crc_out_1_0[22]_net_1 ), .C(feedback_16), .Y(
        \crc_out_1_2[22]_net_1 ));
    AX1C \crc_out_1_3[13]  (.A(N_170_0_0), .B(crc_poly_out_9), .C(
        \crc_out_1_2[13]_net_1 ), .Y(\crc_out_1_3[13]_net_1 ));
    XOR3 \crc_out_1_2[5]  (.A(feedback_1_d0), .B(
        \crc_out_1_0[5]_net_1 ), .C(feedback_0_2), .Y(
        \crc_out_1_2[5]_net_1 ));
    NOR3C \feedback[3]  (.A(crc_poly_size_77), .B(crc_poly_out_3), .C(
        N_170_0), .Y(\feedback_6[3] ));
    XOR3 \crc_out_1_1[18]  (.A(feedback_4_14), .B(crc_in_masked_0_0), 
        .C(feedback_4_15), .Y(crc_out_1_1_14));
    NOR2B \feedback[4]  (.A(crc_poly_out_4), .B(N_170), .Y(
        feedback_5_2));
    XOR3 \crc_out_1_6_RNO_0[9]  (.A(feedback_1_3), .B(\crc_out_1_1[9] )
        , .C(feedback_1_4), .Y(\crc_out_1_3[9] ));
    XOR2 \crc_out_1[9]  (.A(\feedback[9]_net_1 ), .B(
        \crc_out_1_6[9]_net_1 ), .Y(\crc_comb_out[8][9] ));
    NOR2B \feedback[30]  (.A(poly_mux_29), .B(N_170), .Y(
        \feedback[30]_net_1 ));
    XOR2 \crc_out_1[1]  (.A(\feedback[1] ), .B(\crc_comb_out[7]_0 ), 
        .Y(\crc_comb_out[8]_0 ));
    XOR3 \crc_out_1_2[10]  (.A(feedback_3_d0), .B(
        \crc_out_1_0[10]_net_1 ), .C(feedback_4_d0), .Y(
        \crc_out_1_2[10]_net_1 ));
    NOR2B \crc_out_1_6_RNO_2[9]  (.A(crc_init_mux_1), .B(
        crc_poly_size_77), .Y(\un150_crc_init_justified[1] ));
    XOR3 \crc_out_1[29]  (.A(feedback_0_27), .B(
        \crc_out_1_2[29]_net_1 ), .C(\feedback_0[29] ), .Y(
        \crc_comb_out[8]_28 ));
    OR3 \crc_out_1_0_RNINH2GJB2[28]  (.A(un15_crc_out_0), .B(
        crc_out_1_0_0[3]), .C(\un15_crc_out[28] ), .Y(crc_unit_out_0));
    NOR3C \feedback[5]  (.A(crc_poly_size_77), .B(crc_poly_out_5), .C(
        N_170_0), .Y(\feedback_5[5] ));
    AX1C \crc_out_1_0[6]  (.A(N_170_1), .B(poly_mux_0), .C(
        \crc_comb_out[2]_0 ), .Y(\crc_out_1_0[6]_net_1 ));
    NOR2B \feedback[29]  (.A(poly_mux_28), .B(N_170), .Y(
        \feedback_0[29] ));
    XOR3 \crc_out_1_2[19]  (.A(feedback_1_16), .B(
        \crc_out_1_0[19]_net_1 ), .C(feedback_1_17), .Y(
        \crc_out_1_2[19]_net_1 ));
    AX1C \crc_out_1_0[11]  (.A(N_170_0_4), .B(crc_poly_out_4), .C(
        crc_init_mux_3), .Y(\crc_out_1_0[11]_net_1 ));
    AX1C \crc_out_1_1[31]  (.A(N_170_1), .B(poly_mux_25), .C(
        \crc_out_1_0[31]_net_1 ), .Y(\crc_out_1_1[31]_net_1 ));
    XOR3 \crc_out_1[6]  (.A(feedback_6_2), .B(\crc_out_1_3[6]_net_1 ), 
        .C(\feedback_5[6] ), .Y(\crc_comb_out[8]_5 ));
    XOR3 \crc_out_1_2[13]  (.A(feedback_1_6), .B(
        \crc_out_1_0[13]_net_1 ), .C(feedback_2_6), .Y(
        \crc_out_1_2[13]_net_1 ));
    AX1C un2_feedback_6 (.A(N_170_0_2), .B(poly_mux_29), .C(
        un2_feedback_5_net_1), .Y(un2_feedback_6_net_1));
    XOR3 un2_feedback_1 (.A(crc_init_justified[24]), .B(crc_data_in[0])
        , .C(feedback_3_23), .Y(un2_feedback_1_net_1));
    AX1C \crc_out_1_4_RNO_1[15]  (.A(N_170_3), .B(poly_mux_7), .C(
        \un120_crc_init_justified[7] ), .Y(\crc_out_1_0[15] ));
    XOR3 \crc_out_1_6[8]  (.A(feedback_2_4), .B(\crc_out_1_4[8]_net_1 )
        , .C(feedback_4_5), .Y(crc_out_1_6_0));
    XOR3 \crc_out_1_6[11]  (.A(feedback_3_7), .B(
        \crc_out_1_4[11]_net_1 ), .C(feedback_2_8), .Y(crc_out_1_6_3));
    XA1 \crc_out_1_0_RNIOMSNFC2_0[28]  (.A(\feedback_1[28] ), .B(
        \crc_out_1_2[28] ), .C(crc_poly_size_74_0), .Y(
        \un15_crc_out[28] ));
    OR3 \crc_out_1_0_RNIPHJC9N3[28]  (.A(un20_crc_out_16), .B(
        un20_crc_out_0), .C(\un20_crc_out[28] ), .Y(\crc_out_1_1[4] ));
    XA1 \crc_out_1_0_RNIOMSNFC2[28]  (.A(\feedback_1[28] ), .B(
        \crc_out_1_2[28] ), .C(crc_poly_size_77), .Y(crc_unit_out_25));
    NOR3C \feedback[14]  (.A(crc_poly_size_77), .B(crc_poly_out_14), 
        .C(N_170_0), .Y(\feedback_0[14] ));
    AX1 \crc_out_1_0[21]  (.A(crc_poly_size_76_0), .B(
        \crc_comb_out[2]_15 ), .C(feedback_0_15), .Y(
        \crc_out_1_0[21]_net_1 ));
    AX1C un2_feedback_4 (.A(N_170_0_0), .B(poly_mux_27), .C(
        un2_feedback_3_net_1), .Y(un2_feedback_4_net_1));
    XOR3 \crc_out_1_5[23]  (.A(feedback_1_19), .B(
        \crc_out_1_3[23]_net_1 ), .C(feedback_0_20), .Y(
        \crc_out_1_5[23]_net_1 ));
    AX1C \crc_out_1_0_RNICJQ4UA[28]  (.A(N_170_0_2), .B(poly_mux_25), 
        .C(\crc_out_1_0[28]_net_1 ), .Y(\crc_out_1_1[28] ));
    XOR3 \crc_out_1_2[29]  (.A(feedback_25), .B(
        \crc_out_1_0[29]_net_1 ), .C(feedback_26), .Y(
        \crc_out_1_2[29]_net_1 ));
    NOR2B \feedback[26]  (.A(poly_mux_25), .B(N_170), .Y(
        \feedback_1[26] ));
    XOR3 \crc_out_1_4[22]  (.A(feedback_17), .B(
        \crc_out_1_2[22]_net_1 ), .C(feedback_18), .Y(
        \crc_out_1_4[22]_net_1 ));
    XOR3 \crc_out_1_3[20]  (.A(feedback_3_16), .B(
        \crc_out_1_1[20]_net_1 ), .C(feedback_2_17), .Y(crc_out_1_3_14)
        );
    XOR3 \crc_out_1[17]  (.A(feedback_5_14), .B(crc_in_masked_1_0), .C(
        \feedback_5[17] ), .Y(\crc_comb_out[8]_16 ));
    AX1C \crc_out_1_0_RNISA9KP01[28]  (.A(N_170_0_1), .B(poly_mux_26), 
        .C(\crc_out_1_1[28] ), .Y(\crc_out_1_2[28] ));
    AX1C \crc_out_1_0[8]  (.A(N_170_3), .B(poly_mux_0), .C(
        crc_init_mux_0), .Y(\crc_out_1_0[8]_net_1 ));
    AX1C \crc_out_1_0[31]  (.A(N_170_2), .B(poly_mux_24), .C(
        crc_in_masked_0_9), .Y(\crc_out_1_0[31]_net_1 ));
    XOR3 \crc_out_1_5[14]  (.A(feedback_10), .B(
        \crc_out_1_3[14]_net_1 ), .C(feedback_0_11), .Y(
        \crc_out_1_5[14]_net_1 ));
    XOR3 \crc_out_1[7]  (.A(feedback_4_4), .B(\crc_out_1_4[7]_net_1 ), 
        .C(\feedback_6[7] ), .Y(\crc_comb_out[8]_6 ));
    XOR2 \crc_out_1_4[15]  (.A(feedback_11), .B(\crc_out_1_3[15] ), .Y(
        \crc_out_1_4[15]_net_1 ));
    OA1 \feedback[17]  (.A(un84_poly_mux_16), .B(un84_poly_mux_0), .C(
        N_170_0), .Y(\feedback_5[17] ));
    XOR2 un2_feedback_0 (.A(un2_feedback_6_net_1), .B(feedback_30), .Y(
        N_170_0));
    XOR3 \crc_out_1[23]  (.A(feedback_21), .B(\crc_out_1_5[23]_net_1 ), 
        .C(\feedback[23]_net_1 ), .Y(\crc_comb_out[8]_22 ));
    XA1B \crc_in_masked[15]  (.A(feedback_0_14), .B(crc_out_1_5_0[15]), 
        .C(crc_poly_size_76_1), .Y(crc_in_masked_2_0));
    XOR3 \crc_out_1_5[12]  (.A(feedback_2_7), .B(
        \crc_out_1_3[12]_net_1 ), .C(feedback_1_9), .Y(
        \crc_out_1_5[12]_net_1 ));
    XOR3 \crc_out_1_1[14]  (.A(feedback_6_d0), .B(crc_init_mux_6), .C(
        feedback_0_7), .Y(\crc_out_1_1[14]_net_1 ));
    XA1B \crc_in_masked[24]  (.A(feedback_23), .B(crc_in_masked_8), .C(
        crc_poly_size_74_0), .Y(crc_in_masked_3[24]));
    NOR3C \feedback[7]  (.A(crc_poly_size_77), .B(crc_poly_out_7), .C(
        N_170_0), .Y(\feedback_6[7] ));
    XOR2 \crc_out_1_0[28]  (.A(feedback_24), .B(crc_in_masked_9), .Y(
        \crc_out_1_0[28]_net_1 ));
    NOR2B \feedback[28]  (.A(poly_mux_27), .B(N_170), .Y(
        \feedback_1[28] ));
    AX1C \crc_out_1_1[6]  (.A(N_170_5), .B(crc_poly_out_2), .C(
        \crc_out_1_0[6]_net_1 ), .Y(\crc_out_1_1[6]_net_1 ));
    XOR3 \crc_out_1_4_RNO[15]  (.A(feedback_0_9), .B(\crc_out_1_1[15] )
        , .C(feedback_0_10), .Y(\crc_out_1_3[15] ));
    XOR3 \crc_out_1_1[12]  (.A(feedback_2_3), .B(crc_init_mux_4), .C(
        feedback_1_5), .Y(\crc_out_1_1[12]_net_1 ));
    AX1C \crc_out_1_0[3]  (.A(N_170_6), .B(poly_mux_0), .C(
        \crc_comb_out[5] [0]), .Y(\crc_out_1_0[3]_net_1 ));
    AX1C \crc_out_1_0[7]  (.A(N_170_2), .B(poly_mux_0), .C(
        \crc_comb_out[1] [0]), .Y(\crc_out_1_0[7]_net_1 ));
    XOR2 un2_feedback (.A(un2_feedback_6_net_1), .B(feedback_30), .Y(
        N_170));
    XOR3 \crc_out_1_6_RNO_1[9]  (.A(feedback_1_1), .B(
        \un150_crc_init_justified[1] ), .C(feedback_2_1), .Y(
        \crc_out_1_1[9] ));
    XOR2 \crc_out_1_5[15]  (.A(feedback_12), .B(
        \crc_out_1_4[15]_net_1 ), .Y(\crc_out_1_5[15]_net_1 ));
    XOR3 \crc_out_1_2[7]  (.A(feedback_0_1), .B(\crc_out_1_0[7]_net_1 )
        , .C(feedback_1_2), .Y(\crc_out_1_2[7]_net_1 ));
    XOR3 \crc_out_1_4[31]  (.A(feedback_27), .B(
        \crc_out_1_2[31]_net_1 ), .C(feedback_28), .Y(
        \crc_out_1_4[31]_net_1 ));
    XOR3 \crc_out_1_3[23]  (.A(feedback_2_16), .B(
        \crc_out_1_1[23]_net_1 ), .C(feedback_1_18), .Y(
        \crc_out_1_3[23]_net_1 ));
    AX1C \crc_out_1_4_RNO_0[15]  (.A(N_170_2), .B(poly_mux_8), .C(
        \crc_out_1_0[15] ), .Y(\crc_out_1_1[15] ));
    
endmodule


module \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_2 (
       un100_crc_init_justified,
       crc_out_1_2_8,
       un60_crc_init_justified_0,
       un60_crc_init_justified_16,
       un15_crc_init_justified,
       crc_init_justified_1,
       crc_data_in,
       crc_in_masked,
       crc_out_1_1,
       un104_poly_mux_16,
       un104_poly_mux_0,
       un109_poly_mux_16,
       un109_poly_mux_0,
       un79_poly_mux_16,
       un79_poly_mux_0,
       un84_poly_mux_16,
       un84_poly_mux_0,
       un89_poly_mux_16,
       un89_poly_mux_0,
       un94_poly_mux_16,
       un94_poly_mux_0,
       un99_poly_mux_16,
       un99_poly_mux_0,
       feedback_0_18,
       feedback_0_8,
       feedback_0_9,
       feedback_0_7,
       feedback_0_0,
       feedback_0_1,
       feedback_30,
       feedback_12,
       feedback_13,
       feedback_20,
       feedback_21,
       feedback_19,
       feedback_14,
       feedback_24,
       feedback_15,
       feedback_16,
       feedback_17,
       feedback_18,
       feedback_11,
       feedback_5,
       feedback_2,
       feedback_0_d0,
       feedback_4,
       feedback_3,
       feedback_9,
       feedback_10,
       feedback_7,
       feedback_22,
       feedback_6,
       \crc_comb_out[3] ,
       poly_mux_6,
       poly_mux_24,
       poly_mux_23,
       poly_mux_9,
       poly_mux_25,
       poly_mux_19,
       poly_mux_7,
       poly_mux_0,
       poly_mux_17,
       poly_mux_18,
       \crc_comb_out[4]_15 ,
       \crc_comb_out[4]_24 ,
       \crc_comb_out[4]_0 ,
       crc_poly_out_14,
       crc_poly_out_3,
       crc_poly_out_1,
       crc_poly_out_5,
       crc_poly_out_4,
       crc_poly_out_10,
       crc_poly_out_11,
       crc_poly_out_8,
       crc_poly_out_7,
       crc_poly_out_0,
       N_170_0,
       N_170_0_0,
       N_170,
       N_170_1,
       N_170_2,
       crc_poly_size_76_0,
       crc_poly_size_77,
       crc_poly_size_75_0
    );
input  [11:11] un100_crc_init_justified;
output crc_out_1_2_8;
input  un60_crc_init_justified_0;
input  un60_crc_init_justified_16;
input  [28:28] un15_crc_init_justified;
input  [28:28] crc_init_justified_1;
input  [4:4] crc_data_in;
output [15:15] crc_in_masked;
input  [15:15] crc_out_1_1;
input  un104_poly_mux_16;
input  un104_poly_mux_0;
input  un109_poly_mux_16;
input  un109_poly_mux_0;
input  un79_poly_mux_16;
input  un79_poly_mux_0;
input  un84_poly_mux_16;
input  un84_poly_mux_0;
input  un89_poly_mux_16;
input  un89_poly_mux_0;
input  un94_poly_mux_16;
input  un94_poly_mux_0;
input  un99_poly_mux_16;
input  un99_poly_mux_0;
output feedback_0_18;
output feedback_0_8;
output feedback_0_9;
output feedback_0_7;
output feedback_0_0;
output feedback_0_1;
input  feedback_30;
input  feedback_12;
input  feedback_13;
input  feedback_20;
input  feedback_21;
input  feedback_19;
input  feedback_14;
output feedback_24;
output feedback_15;
output feedback_16;
output feedback_17;
output feedback_18;
output feedback_11;
output feedback_5;
output feedback_2;
output feedback_0_d0;
output feedback_4;
output feedback_3;
output feedback_9;
output feedback_10;
output feedback_7;
output feedback_22;
output feedback_6;
input  [23:23] \crc_comb_out[3] ;
input  poly_mux_6;
input  poly_mux_24;
input  poly_mux_23;
input  poly_mux_9;
input  poly_mux_25;
input  poly_mux_19;
input  poly_mux_7;
input  poly_mux_0;
input  poly_mux_17;
input  poly_mux_18;
output \crc_comb_out[4]_15 ;
output \crc_comb_out[4]_24 ;
output \crc_comb_out[4]_0 ;
input  crc_poly_out_14;
input  crc_poly_out_3;
input  crc_poly_out_1;
input  crc_poly_out_5;
input  crc_poly_out_4;
input  crc_poly_out_10;
input  crc_poly_out_11;
input  crc_poly_out_8;
input  crc_poly_out_7;
input  crc_poly_out_0;
output N_170_0;
input  N_170_0_0;
input  N_170;
input  N_170_1;
output N_170_2;
input  crc_poly_size_76_0;
input  crc_poly_size_77;
input  crc_poly_size_75_0;

    wire un2_feedback_2_net_1, \crc_out_1_2[15]_net_1 , 
        \crc_out_1_0[15]_net_1 , \crc_out_1_0[23]_net_1 , 
        un2_feedback_1_net_1, un2_feedback_0_net_1, 
        \feedback[24]_net_1 , GND, VCC;
    
    XOR3 \crc_out_1_2[23]  (.A(feedback_20), .B(
        \crc_out_1_0[23]_net_1 ), .C(feedback_21), .Y(crc_out_1_2_8));
    NOR2B \feedback[10]  (.A(crc_poly_out_10), .B(N_170_2), .Y(
        feedback_9));
    OA1 \feedback[17]  (.A(un84_poly_mux_16), .B(un84_poly_mux_0), .C(
        N_170_0), .Y(feedback_16));
    NOR3C \feedback[5]  (.A(crc_poly_size_77), .B(crc_poly_out_5), .C(
        N_170_2), .Y(feedback_4));
    AX1D \crc_out_1_0[23]  (.A(un60_crc_init_justified_0), .B(
        un60_crc_init_justified_16), .C(feedback_19), .Y(
        \crc_out_1_0[23]_net_1 ));
    NOR3C \feedback[7]  (.A(crc_poly_size_77), .B(crc_poly_out_7), .C(
        N_170_2), .Y(feedback_6));
    VCC VCC_i (.Y(VCC));
    XOR3 \crc_out_1_2[15]  (.A(feedback_12), .B(
        \crc_out_1_0[15]_net_1 ), .C(feedback_13), .Y(
        \crc_out_1_2[15]_net_1 ));
    AX1C \crc_out_1[15]  (.A(N_170_0), .B(poly_mux_9), .C(
        \crc_out_1_2[15]_net_1 ), .Y(\crc_comb_out[4]_15 ));
    NOR2B \feedback[23]  (.A(poly_mux_17), .B(N_170_2), .Y(feedback_22)
        );
    AX1C un2_feedback_1 (.A(N_170_1), .B(poly_mux_23), .C(
        un2_feedback_0_net_1), .Y(un2_feedback_1_net_1));
    NOR2B \feedback[8]  (.A(crc_poly_out_8), .B(N_170_2), .Y(
        feedback_7));
    AX1D un2_feedback_0 (.A(un15_crc_init_justified[28]), .B(
        crc_init_justified_1[28]), .C(crc_data_in[4]), .Y(
        un2_feedback_0_net_1));
    NOR3C \feedback[14]  (.A(crc_poly_size_77), .B(crc_poly_out_14), 
        .C(N_170_0), .Y(feedback_0_1));
    AX1C \crc_out_1_0[15]  (.A(N_170_0_0), .B(poly_mux_6), .C(
        un100_crc_init_justified[11]), .Y(\crc_out_1_0[15]_net_1 ));
    NOR2B \feedback[12]  (.A(poly_mux_6), .B(N_170_2), .Y(feedback_11));
    OA1 \feedback[21]  (.A(un104_poly_mux_16), .B(un104_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_8));
    OA1 \feedback[19]  (.A(un94_poly_mux_16), .B(un94_poly_mux_0), .C(
        N_170_0), .Y(feedback_18));
    XOR2 un2_feedback_0_0 (.A(un2_feedback_2_net_1), .B(feedback_30), 
        .Y(N_170_0));
    NOR2B \feedback[25]  (.A(poly_mux_19), .B(N_170_2), .Y(feedback_24)
        );
    AX1C un2_feedback_2 (.A(N_170), .B(poly_mux_24), .C(
        un2_feedback_1_net_1), .Y(un2_feedback_2_net_1));
    OA1 \feedback[20]  (.A(un99_poly_mux_16), .B(un99_poly_mux_0), .C(
        N_170_0), .Y(feedback_0_7));
    AX1 \crc_out_1[24]  (.A(crc_poly_size_75_0), .B(
        \crc_comb_out[3] [23]), .C(\feedback[24]_net_1 ), .Y(
        \crc_comb_out[4]_24 ));
    XOR2 un2_feedback (.A(un2_feedback_2_net_1), .B(feedback_30), .Y(
        N_170_2));
    NOR2B \feedback[6]  (.A(poly_mux_0), .B(N_170_2), .Y(feedback_5));
    GND GND_i (.Y(GND));
    NOR2B \feedback[31]  (.A(poly_mux_25), .B(N_170_2), .Y(
        feedback_0_18));
    NOR2B \feedback[24]  (.A(poly_mux_18), .B(N_170_2), .Y(
        \feedback[24]_net_1 ));
    OA1 \feedback[22]  (.A(un109_poly_mux_16), .B(un109_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_9));
    NOR2B \feedback[0]  (.A(crc_poly_out_0), .B(N_170_2), .Y(
        \crc_comb_out[4]_0 ));
    XA1B \crc_in_masked[15]  (.A(feedback_14), .B(crc_out_1_1[15]), .C(
        crc_poly_size_76_0), .Y(crc_in_masked[15]));
    NOR2B \feedback[4]  (.A(crc_poly_out_4), .B(N_170_2), .Y(
        feedback_3));
    NOR2B \feedback[13]  (.A(poly_mux_7), .B(N_170_2), .Y(feedback_0_0)
        );
    NOR2B \feedback[1]  (.A(crc_poly_out_1), .B(N_170_2), .Y(
        feedback_0_d0));
    NOR2B \feedback[3]  (.A(crc_poly_out_3), .B(N_170_2), .Y(
        feedback_2));
    OA1 \feedback[18]  (.A(un89_poly_mux_16), .B(un89_poly_mux_0), .C(
        N_170_0), .Y(feedback_17));
    OA1 \feedback[16]  (.A(un79_poly_mux_16), .B(un79_poly_mux_0), .C(
        N_170_0), .Y(feedback_15));
    NOR3C \feedback[11]  (.A(crc_poly_size_77), .B(crc_poly_out_11), 
        .C(N_170_0), .Y(feedback_10));
    
endmodule


module \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_5 (
       crc_out_1_5,
       un115_crc_init_justified,
       un75_crc_init_justified_16,
       un75_crc_init_justified_0,
       un30_crc_init_justified,
       crc_init_justified_1,
       crc_data_in,
       \crc_comb_out[7]_0 ,
       \crc_comb_out[7]_23 ,
       crc_out_1_4_0,
       un104_poly_mux_16,
       un104_poly_mux_0,
       un109_poly_mux_16,
       un109_poly_mux_0,
       un84_poly_mux_16,
       un84_poly_mux_0,
       un94_poly_mux_16,
       un94_poly_mux_0,
       un99_poly_mux_16,
       un99_poly_mux_0,
       un79_poly_mux_16,
       un79_poly_mux_0,
       crc_in_masked_8,
       crc_in_masked_0,
       crc_out_1_4_0_d0,
       un89_poly_mux_16,
       un89_poly_mux_0,
       feedback_0_14,
       feedback_0_22,
       feedback_0_12,
       feedback_0_13,
       feedback_0_8,
       feedback_0_10,
       feedback_0_11,
       feedback_0_5,
       feedback_0_0,
       feedback_0_3,
       feedback_0_4,
       feedback_0_6,
       feedback_0_2,
       feedback_0_9,
       feedback_0_1,
       poly_mux_29,
       poly_mux_28,
       poly_mux_27,
       poly_mux_26,
       poly_mux_25,
       poly_mux_30,
       poly_mux_23,
       poly_mux_24,
       poly_mux_14,
       poly_mux_7,
       poly_mux_8,
       poly_mux_0,
       poly_mux_5,
       poly_mux_11,
       poly_mux_22,
       poly_mux_12,
       poly_mux_9,
       feedback_30,
       feedback_12,
       feedback_13,
       feedback_10,
       feedback_11,
       feedback_8,
       feedback_9,
       feedback_19,
       feedback_20,
       feedback_17,
       feedback_18,
       feedback_16,
       feedback_21,
       feedback_25,
       feedback_27,
       feedback_29,
       feedback_23,
       feedback_24,
       feedback_14,
       feedback_7,
       feedback_0_d0,
       feedback_5,
       feedback_3,
       feedback_4,
       feedback_6,
       feedback_15,
       feedback_1,
       feedback_2,
       crc_poly_out_0,
       crc_poly_out_14,
       crc_poly_out_4,
       crc_poly_out_5,
       crc_poly_out_7,
       crc_poly_out_11,
       crc_poly_out_2,
       crc_poly_out_3,
       N_170_0,
       N_170,
       N_170_0_0,
       N_170_1,
       N_170_2,
       N_170_3,
       crc_poly_size_75_0,
       crc_poly_size_77,
       crc_poly_size_76_0
    );
output [15:15] crc_out_1_5;
input  [8:8] un115_crc_init_justified;
input  un75_crc_init_justified_16;
input  un75_crc_init_justified_0;
input  [25:25] un30_crc_init_justified;
input  [25:25] crc_init_justified_1;
input  [1:1] crc_data_in;
output \crc_comb_out[7]_0 ;
output \crc_comb_out[7]_23 ;
input  [23:23] crc_out_1_4_0;
input  un104_poly_mux_16;
input  un104_poly_mux_0;
input  un109_poly_mux_16;
input  un109_poly_mux_0;
input  un84_poly_mux_16;
input  un84_poly_mux_0;
input  un94_poly_mux_16;
input  un94_poly_mux_0;
input  un99_poly_mux_16;
input  un99_poly_mux_0;
input  un79_poly_mux_16;
input  un79_poly_mux_0;
output crc_in_masked_8;
output crc_in_masked_0;
input  crc_out_1_4_0_d0;
input  un89_poly_mux_16;
input  un89_poly_mux_0;
input  feedback_0_14;
output feedback_0_22;
output feedback_0_12;
output feedback_0_13;
output feedback_0_8;
output feedback_0_10;
output feedback_0_11;
output feedback_0_5;
output feedback_0_0;
output feedback_0_3;
output feedback_0_4;
input  feedback_0_6;
output feedback_0_2;
output feedback_0_9;
output feedback_0_1;
input  poly_mux_29;
input  poly_mux_28;
input  poly_mux_27;
input  poly_mux_26;
input  poly_mux_25;
input  poly_mux_30;
input  poly_mux_23;
input  poly_mux_24;
input  poly_mux_14;
input  poly_mux_7;
input  poly_mux_8;
input  poly_mux_0;
input  poly_mux_5;
input  poly_mux_11;
input  poly_mux_22;
input  poly_mux_12;
input  poly_mux_9;
input  feedback_30;
input  feedback_12;
input  feedback_13;
input  feedback_10;
input  feedback_11;
input  feedback_8;
input  feedback_9;
input  feedback_19;
input  feedback_20;
input  feedback_17;
input  feedback_18;
input  feedback_16;
input  feedback_21;
output feedback_25;
output feedback_27;
output feedback_29;
output feedback_23;
output feedback_24;
output feedback_14;
output feedback_7;
output feedback_0_d0;
output feedback_5;
output feedback_3;
output feedback_4;
output feedback_6;
output feedback_15;
output feedback_1;
output feedback_2;
input  crc_poly_out_0;
input  crc_poly_out_14;
input  crc_poly_out_4;
input  crc_poly_out_5;
input  crc_poly_out_7;
input  crc_poly_out_11;
input  crc_poly_out_2;
input  crc_poly_out_3;
output N_170_0;
input  N_170;
input  N_170_0_0;
input  N_170_1;
input  N_170_2;
input  N_170_3;
input  crc_poly_size_75_0;
input  crc_poly_size_77;
input  crc_poly_size_76_0;

    wire un2_feedback_5_net_1, \crc_out_1_3[15]_net_1 , 
        \crc_out_1_1[15]_net_1 , \crc_out_1_4[23]_net_1 , 
        \crc_out_1_2[23]_net_1 , \crc_out_1_0[23]_net_1 , 
        un2_feedback_4_net_1, un2_feedback_3_net_1, 
        un2_feedback_2_net_1, un2_feedback_1_net_1, 
        un2_feedback_0_net_1, N_170_4, \feedback[23]_net_1 , GND, VCC;
    
    NOR2B \feedback[15]  (.A(poly_mux_14), .B(N_170_4), .Y(feedback_14)
        );
    XOR3 \crc_out_1_2[23]  (.A(feedback_17), .B(
        \crc_out_1_0[23]_net_1 ), .C(feedback_18), .Y(
        \crc_out_1_2[23]_net_1 ));
    NOR2B \feedback[10]  (.A(poly_mux_9), .B(N_170_4), .Y(feedback_0_1)
        );
    XOR3 \crc_out_1_4[23]  (.A(feedback_19), .B(
        \crc_out_1_2[23]_net_1 ), .C(feedback_20), .Y(
        \crc_out_1_4[23]_net_1 ));
    OA1 \feedback[17]  (.A(un84_poly_mux_16), .B(un84_poly_mux_0), .C(
        N_170_0), .Y(feedback_0_8));
    XOR3 \crc_out_1_3[15]  (.A(feedback_10), .B(
        \crc_out_1_1[15]_net_1 ), .C(feedback_11), .Y(
        \crc_out_1_3[15]_net_1 ));
    NOR2B \feedback[5]  (.A(crc_poly_out_5), .B(N_170_4), .Y(
        feedback_4));
    XA1B \crc_in_masked[23]  (.A(feedback_0_14), .B(crc_out_1_4_0[23]), 
        .C(crc_poly_size_75_0), .Y(crc_in_masked_8));
    AX1D \crc_out_1_0[23]  (.A(un75_crc_init_justified_16), .B(
        un75_crc_init_justified_0), .C(feedback_16), .Y(
        \crc_out_1_0[23]_net_1 ));
    NOR3C \feedback[7]  (.A(crc_poly_size_77), .B(crc_poly_out_7), .C(
        N_170_0), .Y(feedback_6));
    VCC VCC_i (.Y(VCC));
    NOR2B \feedback[23]  (.A(poly_mux_22), .B(N_170_4), .Y(
        \feedback[23]_net_1 ));
    AX1C un2_feedback_1 (.A(N_170_3), .B(poly_mux_25), .C(
        un2_feedback_0_net_1), .Y(un2_feedback_1_net_1));
    NOR2B \feedback[8]  (.A(poly_mux_7), .B(N_170_4), .Y(feedback_7));
    AX1D un2_feedback_0 (.A(un30_crc_init_justified[25]), .B(
        crc_init_justified_1[25]), .C(crc_data_in[1]), .Y(
        un2_feedback_0_net_1));
    NOR2B \feedback[28]  (.A(poly_mux_27), .B(N_170_4), .Y(feedback_27)
        );
    NOR3C \feedback[14]  (.A(crc_poly_size_77), .B(crc_poly_out_14), 
        .C(N_170_0), .Y(feedback_0_5));
    NOR2B \feedback[26]  (.A(poly_mux_25), .B(N_170_4), .Y(feedback_25)
        );
    NOR2B \feedback[12]  (.A(poly_mux_11), .B(N_170_4), .Y(
        feedback_0_3));
    NOR3C \feedback[2]  (.A(crc_poly_size_77), .B(crc_poly_out_2), .C(
        N_170_0), .Y(feedback_1));
    OA1 \feedback[21]  (.A(un104_poly_mux_16), .B(un104_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_12));
    OA1 \feedback[19]  (.A(un94_poly_mux_16), .B(un94_poly_mux_0), .C(
        N_170_0), .Y(feedback_0_10));
    XOR2 un2_feedback_0_0 (.A(un2_feedback_5_net_1), .B(feedback_30), 
        .Y(N_170_0));
    NOR2B \feedback[25]  (.A(poly_mux_24), .B(N_170_4), .Y(feedback_24)
        );
    NOR2B \feedback[9]  (.A(poly_mux_8), .B(N_170_4), .Y(feedback_0_0));
    AX1C un2_feedback_2 (.A(N_170_2), .B(poly_mux_26), .C(
        un2_feedback_1_net_1), .Y(un2_feedback_2_net_1));
    OA1 \feedback[20]  (.A(un99_poly_mux_16), .B(un99_poly_mux_0), .C(
        N_170_0), .Y(feedback_0_11));
    XOR2 un2_feedback (.A(un2_feedback_5_net_1), .B(feedback_30), .Y(
        N_170_4));
    NOR2B \feedback[6]  (.A(poly_mux_5), .B(N_170_4), .Y(feedback_5));
    GND GND_i (.Y(GND));
    AX1C un2_feedback_5 (.A(N_170), .B(poly_mux_29), .C(
        un2_feedback_4_net_1), .Y(un2_feedback_5_net_1));
    AX1C un2_feedback_4 (.A(N_170_0_0), .B(poly_mux_28), .C(
        un2_feedback_3_net_1), .Y(un2_feedback_4_net_1));
    NOR2B \feedback[31]  (.A(poly_mux_30), .B(N_170_4), .Y(
        feedback_0_22));
    AX1C un2_feedback_3 (.A(N_170_1), .B(poly_mux_27), .C(
        un2_feedback_2_net_1), .Y(un2_feedback_3_net_1));
    NOR2B \feedback[24]  (.A(poly_mux_23), .B(N_170_4), .Y(feedback_23)
        );
    NOR2B \feedback[30]  (.A(poly_mux_29), .B(N_170_4), .Y(feedback_29)
        );
    OA1 \feedback[22]  (.A(un109_poly_mux_16), .B(un109_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_13));
    XOR3 \crc_out_1[23]  (.A(feedback_21), .B(\crc_out_1_4[23]_net_1 ), 
        .C(\feedback[23]_net_1 ), .Y(\crc_comb_out[7]_23 ));
    XOR3 \crc_out_1_5[15]  (.A(feedback_12), .B(
        \crc_out_1_3[15]_net_1 ), .C(feedback_13), .Y(crc_out_1_5[15]));
    AND2 \feedback[0]  (.A(N_170_0), .B(crc_poly_out_0), .Y(
        \crc_comb_out[7]_0 ));
    XA1B \crc_in_masked[15]  (.A(feedback_0_6), .B(crc_out_1_4_0_d0), 
        .C(crc_poly_size_76_0), .Y(crc_in_masked_0));
    NOR3C \feedback[4]  (.A(crc_poly_size_77), .B(crc_poly_out_4), .C(
        N_170_0), .Y(feedback_3));
    NOR2B \feedback[13]  (.A(poly_mux_12), .B(N_170_4), .Y(
        feedback_0_4));
    NOR2B \feedback[1]  (.A(poly_mux_0), .B(N_170_4), .Y(feedback_0_d0)
        );
    NOR3C \feedback[3]  (.A(crc_poly_size_77), .B(crc_poly_out_3), .C(
        N_170_0), .Y(feedback_2));
    OA1 \feedback[18]  (.A(un89_poly_mux_16), .B(un89_poly_mux_0), .C(
        N_170_0), .Y(feedback_0_9));
    OA1 \feedback[16]  (.A(un79_poly_mux_16), .B(un79_poly_mux_0), .C(
        N_170_0), .Y(feedback_15));
    XOR3 \crc_out_1_1[15]  (.A(feedback_8), .B(
        un115_crc_init_justified[8]), .C(feedback_9), .Y(
        \crc_out_1_1[15]_net_1 ));
    NOR3C \feedback[11]  (.A(crc_poly_size_77), .B(crc_poly_out_11), 
        .C(N_170_0), .Y(feedback_0_2));
    
endmodule


module \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_1 (
       \crc_comb_out[2] ,
       crc_out_1_1,
       un95_crc_init_justified,
       un55_crc_init_justified_16,
       un55_crc_init_justified_0,
       un10_crc_init_justified,
       crc_init_justified_1,
       crc_data_in,
       \crc_comb_out[3] ,
       crc_in_masked_1,
       crc_out_1_0_1,
       un104_poly_mux_16,
       un104_poly_mux_0,
       un79_poly_mux_16,
       un79_poly_mux_0,
       un84_poly_mux_16,
       un84_poly_mux_0,
       un89_poly_mux_16,
       un89_poly_mux_0,
       un94_poly_mux_16,
       un94_poly_mux_0,
       un99_poly_mux_16,
       un99_poly_mux_0,
       crc_poly_out_9,
       crc_poly_out_3,
       crc_poly_out_0,
       crc_poly_out_2,
       crc_poly_out_1,
       crc_poly_out_5,
       crc_poly_out_12,
       feedback_0_11,
       feedback_0_18,
       feedback_0_8,
       feedback_0_0,
       feedback_0_1,
       feedback_0_9,
       un109_poly_mux_16,
       un109_poly_mux_0,
       feedback_29,
       feedback_11,
       feedback_12,
       feedback_19,
       feedback_20,
       feedback_14,
       feedback_15,
       feedback_16,
       feedback_17,
       feedback_18,
       feedback_9,
       feedback_10,
       feedback_13,
       feedback_6,
       feedback_3,
       feedback_0_d0,
       feedback_2,
       feedback_1,
       feedback_7,
       feedback_8,
       feedback_5,
       feedback_4,
       poly_mux_18,
       poly_mux_24,
       poly_mux_25,
       poly_mux_6,
       poly_mux_7,
       poly_mux_9,
       poly_mux_2,
       poly_mux_3,
       poly_mux_4,
       poly_mux_0,
       poly_mux_17,
       N_170_0,
       crc_poly_size_75,
       N_170,
       N_170_0_0,
       crc_poly_size_74_0,
       crc_poly_size_77
    );
input  [23:23] \crc_comb_out[2] ;
output [15:15] crc_out_1_1;
input  [12:12] un95_crc_init_justified;
input  un55_crc_init_justified_16;
input  un55_crc_init_justified_0;
input  [29:29] un10_crc_init_justified;
input  [29:29] crc_init_justified_1;
input  [5:5] crc_data_in;
output [24:23] \crc_comb_out[3] ;
output crc_in_masked_1;
input  crc_out_1_0_1;
input  un104_poly_mux_16;
input  un104_poly_mux_0;
input  un79_poly_mux_16;
input  un79_poly_mux_0;
input  un84_poly_mux_16;
input  un84_poly_mux_0;
input  un89_poly_mux_16;
input  un89_poly_mux_0;
input  un94_poly_mux_16;
input  un94_poly_mux_0;
input  un99_poly_mux_16;
input  un99_poly_mux_0;
input  crc_poly_out_9;
input  crc_poly_out_3;
input  crc_poly_out_0;
input  crc_poly_out_2;
input  crc_poly_out_1;
input  crc_poly_out_5;
input  crc_poly_out_12;
input  feedback_0_11;
output feedback_0_18;
output feedback_0_8;
output feedback_0_0;
output feedback_0_1;
output feedback_0_9;
input  un109_poly_mux_16;
input  un109_poly_mux_0;
input  feedback_29;
input  feedback_11;
input  feedback_12;
input  feedback_19;
input  feedback_20;
output feedback_14;
output feedback_15;
output feedback_16;
output feedback_17;
output feedback_18;
output feedback_9;
output feedback_10;
output feedback_13;
output feedback_6;
output feedback_3;
output feedback_0_d0;
output feedback_2;
output feedback_1;
output feedback_7;
output feedback_8;
output feedback_5;
output feedback_4;
input  poly_mux_18;
input  poly_mux_24;
input  poly_mux_25;
input  poly_mux_6;
input  poly_mux_7;
input  poly_mux_9;
input  poly_mux_2;
input  poly_mux_3;
input  poly_mux_4;
input  poly_mux_0;
input  poly_mux_17;
output N_170_0;
input  crc_poly_size_75;
output N_170;
input  N_170_0_0;
input  crc_poly_size_74_0;
input  crc_poly_size_77;

    wire un2_feedback_1_net_1, \crc_in_masked[23]_net_1 , 
        \feedback[24]_net_1 , \crc_out_1_0[23]_net_1 , 
        un2_feedback_0_net_1, \feedback[23]_net_1 , GND, VCC;
    
    NOR2B \feedback[15]  (.A(poly_mux_9), .B(N_170), .Y(feedback_13));
    NOR2B \feedback[10]  (.A(poly_mux_4), .B(N_170), .Y(feedback_8));
    OA1 \feedback[17]  (.A(un84_poly_mux_16), .B(un84_poly_mux_0), .C(
        N_170_0), .Y(feedback_15));
    NOR3C \feedback[5]  (.A(crc_poly_size_77), .B(crc_poly_out_3), .C(
        N_170_0), .Y(feedback_3));
    NOR2A \crc_in_masked[23]  (.A(\crc_comb_out[2] [23]), .B(
        crc_poly_size_75), .Y(\crc_in_masked[23]_net_1 ));
    AX1D \crc_out_1_0[23]  (.A(un55_crc_init_justified_16), .B(
        un55_crc_init_justified_0), .C(feedback_19), .Y(
        \crc_out_1_0[23]_net_1 ));
    NOR3C \feedback[7]  (.A(crc_poly_size_77), .B(crc_poly_out_5), .C(
        N_170_0), .Y(feedback_5));
    VCC VCC_i (.Y(VCC));
    NOR2B \feedback[23]  (.A(poly_mux_17), .B(N_170), .Y(
        \feedback[23]_net_1 ));
    AX1C un2_feedback_1 (.A(N_170_0_0), .B(poly_mux_24), .C(
        un2_feedback_0_net_1), .Y(un2_feedback_1_net_1));
    NOR2B \feedback[8]  (.A(poly_mux_2), .B(N_170), .Y(feedback_6));
    AX1D un2_feedback_0 (.A(un10_crc_init_justified[29]), .B(
        crc_init_justified_1[29]), .C(crc_data_in[5]), .Y(
        un2_feedback_0_net_1));
    NOR3C \feedback[14]  (.A(crc_poly_size_77), .B(crc_poly_out_12), 
        .C(N_170_0), .Y(feedback_0_1));
    NOR2B \feedback[12]  (.A(poly_mux_6), .B(N_170), .Y(feedback_10));
    NOR3C \feedback[2]  (.A(crc_poly_size_77), .B(crc_poly_out_0), .C(
        N_170_0), .Y(feedback_0_d0));
    OA1 \feedback[21]  (.A(un104_poly_mux_16), .B(un104_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_8));
    OA1 \feedback[19]  (.A(un94_poly_mux_16), .B(un94_poly_mux_0), .C(
        N_170_0), .Y(feedback_17));
    XA1B \crc_in_masked[24]  (.A(feedback_0_11), .B(crc_out_1_0_1), .C(
        crc_poly_size_74_0), .Y(crc_in_masked_1));
    XOR2 un2_feedback_0_0 (.A(un2_feedback_1_net_1), .B(feedback_29), 
        .Y(N_170_0));
    NOR2B \feedback[9]  (.A(poly_mux_3), .B(N_170), .Y(feedback_7));
    OA1 \feedback[20]  (.A(un99_poly_mux_16), .B(un99_poly_mux_0), .C(
        N_170_0), .Y(feedback_18));
    XOR2 \crc_out_1[24]  (.A(\feedback[24]_net_1 ), .B(
        \crc_in_masked[23]_net_1 ), .Y(\crc_comb_out[3] [24]));
    XOR2 un2_feedback (.A(un2_feedback_1_net_1), .B(feedback_29), .Y(
        N_170));
    NOR2B \feedback[6]  (.A(poly_mux_0), .B(N_170), .Y(feedback_4));
    GND GND_i (.Y(GND));
    NOR2B \feedback[31]  (.A(poly_mux_25), .B(N_170), .Y(feedback_0_18)
        );
    AND2 \feedback[24]  (.A(N_170), .B(poly_mux_18), .Y(
        \feedback[24]_net_1 ));
    OA1 \feedback[22]  (.A(un109_poly_mux_16), .B(un109_poly_mux_0), 
        .C(N_170_0), .Y(feedback_0_9));
    XOR3 \crc_out_1[23]  (.A(feedback_20), .B(\crc_out_1_0[23]_net_1 ), 
        .C(\feedback[23]_net_1 ), .Y(\crc_comb_out[3] [23]));
    NOR3C \feedback[4]  (.A(crc_poly_size_77), .B(crc_poly_out_2), .C(
        N_170_0), .Y(feedback_2));
    NOR2B \feedback[13]  (.A(poly_mux_7), .B(N_170), .Y(feedback_0_0));
    NOR3C \feedback[3]  (.A(crc_poly_size_77), .B(crc_poly_out_1), .C(
        N_170_0), .Y(feedback_1));
    OA1 \feedback[18]  (.A(un89_poly_mux_16), .B(un89_poly_mux_0), .C(
        N_170_0), .Y(feedback_16));
    OA1 \feedback[16]  (.A(un79_poly_mux_16), .B(un79_poly_mux_0), .C(
        N_170_0), .Y(feedback_14));
    XOR3 \crc_out_1_1[15]  (.A(feedback_11), .B(
        un95_crc_init_justified[12]), .C(feedback_12), .Y(
        crc_out_1_1[15]));
    NOR3C \feedback[11]  (.A(crc_poly_size_77), .B(crc_poly_out_9), .C(
        N_170_0), .Y(feedback_9));
    
endmodule


module \crc_comb_32s_4294967295_genblk4[0].CRC_COMB (
       crc_data_in,
       crc_init_justified,
       un79_poly_mux_16,
       un79_poly_mux_0,
       un84_poly_mux_16,
       un84_poly_mux_0,
       un89_poly_mux_16,
       un89_poly_mux_0,
       un94_poly_mux_16,
       un94_poly_mux_0,
       un109_poly_mux_16,
       un109_poly_mux_0,
       un99_poly_mux_16,
       un99_poly_mux_0,
       \crc_comb_out[1] ,
       crc_poly_out_14,
       crc_poly_out_3,
       crc_poly_out_11,
       crc_poly_out_0,
       crc_poly_out_2,
       crc_poly_out_7,
       crc_poly_out_5,
       poly_mux_4,
       poly_mux_16,
       poly_mux_15,
       poly_mux_22,
       poly_mux_0,
       feedback_11,
       feedback_12,
       feedback_23,
       feedback_14,
       feedback_15,
       feedback_22,
       feedback_1,
       feedback_16,
       feedback_17,
       feedback_20,
       feedback_9,
       feedback_18,
       feedback_0,
       feedback_5,
       feedback_29,
       feedback_3,
       feedback_7,
       feedback_19,
       un104_poly_mux_16,
       un104_poly_mux_0,
       N_170_0,
       N_170,
       crc_poly_size_77
    );
input  [7:7] crc_data_in;
input  [31:31] crc_init_justified;
input  un79_poly_mux_16;
input  un79_poly_mux_0;
input  un84_poly_mux_16;
input  un84_poly_mux_0;
input  un89_poly_mux_16;
input  un89_poly_mux_0;
input  un94_poly_mux_16;
input  un94_poly_mux_0;
input  un109_poly_mux_16;
input  un109_poly_mux_0;
input  un99_poly_mux_16;
input  un99_poly_mux_0;
output [0:0] \crc_comb_out[1] ;
input  crc_poly_out_14;
input  crc_poly_out_3;
input  crc_poly_out_11;
input  crc_poly_out_0;
input  crc_poly_out_2;
input  crc_poly_out_7;
input  crc_poly_out_5;
input  poly_mux_4;
input  poly_mux_16;
input  poly_mux_15;
input  poly_mux_22;
input  poly_mux_0;
output feedback_11;
output feedback_12;
output feedback_23;
output feedback_14;
output feedback_15;
output feedback_22;
output feedback_1;
output feedback_16;
output feedback_17;
output feedback_20;
output feedback_9;
output feedback_18;
output feedback_0;
output feedback_5;
output feedback_29;
output feedback_3;
output feedback_7;
output feedback_19;
input  un104_poly_mux_16;
input  un104_poly_mux_0;
output N_170_0;
output N_170;
input  crc_poly_size_77;

    wire GND, VCC;
    
    NOR3C \feedback[2]  (.A(crc_poly_size_77), .B(crc_poly_out_2), .C(
        N_170), .Y(feedback_0));
    OA1 \feedback[16]  (.A(un79_poly_mux_16), .B(un79_poly_mux_0), .C(
        N_170_0), .Y(feedback_14));
    NOR3C \feedback[7]  (.A(crc_poly_size_77), .B(crc_poly_out_7), .C(
        N_170), .Y(feedback_5));
    OA1 \feedback[17]  (.A(un84_poly_mux_16), .B(un84_poly_mux_0), .C(
        N_170_0), .Y(feedback_15));
    NOR2B \feedback[13]  (.A(poly_mux_4), .B(N_170), .Y(feedback_11));
    XOR2 un2_feedback_0 (.A(crc_data_in[7]), .B(crc_init_justified[31])
        , .Y(N_170_0));
    OA1 \feedback[22]  (.A(un109_poly_mux_16), .B(un109_poly_mux_0), 
        .C(N_170_0), .Y(feedback_20));
    VCC VCC_i (.Y(VCC));
    OA1 \feedback[19]  (.A(un94_poly_mux_16), .B(un94_poly_mux_0), .C(
        N_170_0), .Y(feedback_17));
    OA1 \feedback[21]  (.A(un104_poly_mux_16), .B(un104_poly_mux_0), 
        .C(N_170_0), .Y(feedback_19));
    NOR2B \feedback[0]  (.A(crc_poly_out_0), .B(N_170), .Y(
        \crc_comb_out[1] [0]));
    GND GND_i (.Y(GND));
    NOR3C \feedback[11]  (.A(crc_poly_size_77), .B(crc_poly_out_11), 
        .C(N_170_0), .Y(feedback_9));
    NOR2B \feedback[24]  (.A(poly_mux_15), .B(N_170), .Y(feedback_22));
    NOR2B \feedback[9]  (.A(poly_mux_0), .B(N_170), .Y(feedback_7));
    OA1 \feedback[18]  (.A(un89_poly_mux_16), .B(un89_poly_mux_0), .C(
        N_170_0), .Y(feedback_16));
    NOR3C \feedback[14]  (.A(crc_poly_size_77), .B(crc_poly_out_14), 
        .C(N_170_0), .Y(feedback_12));
    NOR3C \feedback[5]  (.A(crc_poly_size_77), .B(crc_poly_out_5), .C(
        N_170), .Y(feedback_3));
    OA1 \feedback[20]  (.A(un99_poly_mux_16), .B(un99_poly_mux_0), .C(
        N_170_0), .Y(feedback_18));
    XOR2 un2_feedback (.A(crc_data_in[7]), .B(crc_init_justified[31]), 
        .Y(N_170));
    NOR3C \feedback[3]  (.A(crc_poly_size_77), .B(crc_poly_out_3), .C(
        N_170), .Y(feedback_1));
    NOR2B \feedback[31]  (.A(poly_mux_22), .B(N_170), .Y(feedback_29));
    NOR2B \feedback[25]  (.A(poly_mux_16), .B(N_170), .Y(feedback_23));
    
endmodule


module crc_parallel_32s_8s_4294967295_0(
       crc_poly_out,
       crc_init_mux,
       crc_data_in,
       crc_unit_out,
       crc_poly_size_76,
       crc_poly_size_77,
       crc_poly_size_74,
       crc_poly_size_75_0,
       crc_poly_size_76_0,
       crc_poly_size_74_0,
       crc_poly_size_76_1,
       crc_poly_size_75
    );
input  [31:0] crc_poly_out;
input  [31:0] crc_init_mux;
input  [7:0] crc_data_in;
output [31:0] crc_unit_out;
input  crc_poly_size_76;
input  crc_poly_size_77;
input  crc_poly_size_74;
input  crc_poly_size_75_0;
input  crc_poly_size_76_0;
input  crc_poly_size_74_0;
input  crc_poly_size_76_1;
input  crc_poly_size_75;

    wire \un20_crc_init_justified[11]_net_1 , 
        \un15_crc_init_justified[12]_net_1 , \un5_crc_out[1]_net_1 , 
        \crc_comb_out[8][1] , \un5_crc_out[26]_net_1 , 
        \crc_comb_out[8][26] , \un75_crc_out[15]_net_1 , 
        \crc_comb_out[8][15] , \un75_crc_out[31] , 
        \crc_out_1_1[1]_net_1 , \un5_crc_out[25] , \crc_out_1_0[1] , 
        \crc_init_justified_1[28]_net_1 , 
        \crc_init_justified_0[28]_net_1 , \un15_crc_init_justified[4] , 
        \un15_crc_init_justified[3] , \crc_init_justified_1[27]_net_1 , 
        \crc_init_justified_0[27]_net_1 , \un20_crc_init_justified[3] , 
        \un20_crc_init_justified[2] , \crc_out_1_1[5]_net_1 , 
        \crc_comb_out[8][29] , \crc_out_1_0[5]_net_1 , 
        \crc_comb_out[8][5] , \un25_crc_out[21]_net_1 , 
        \crc_out_1_0[6]_net_1 , \crc_comb_out[8][6] , 
        \un30_crc_out[22]_net_1 , \crc_out_1_0[2]_net_1 , 
        \crc_comb_out[8][2] , \un10_crc_out[18]_net_1 , 
        \crc_comb_out[8][17] , \crc_out_1_0[3]_net_1 , 
        \crc_comb_out[8][3] , \un15_crc_out[19]_net_1 , 
        \crc_out_1_0[7]_net_1 , \crc_comb_out[8][23] , 
        \un35_crc_out[7]_net_1 , \crc_out_1_0[0]_net_1 , 
        \un1_crc_out_0[0] , N_170_0, \un1_crc_out[24] , 
        \poly_mux_0[31]_net_1 , \un154_poly_mux[6] , 
        \poly_mux_0[29]_net_1 , \un144_poly_mux[5]_net_1 , 
        \poly_mux_0[27]_net_1 , \un134_poly_mux[3]_net_1 , 
        \poly_mux_1[25]_net_1 , \un124_poly_mux[1]_net_1 , 
        \un124_poly_mux[0]_net_1 , \un124_poly_mux[9]_net_1 , 
        \poly_mux_1[30]_net_1 , \un149_poly_mux[6]_net_1 , 
        \un149_poly_mux[5]_net_1 , \un149_poly_mux[14]_net_1 , 
        \poly_mux_1[28]_net_1 , \un139_poly_mux[4]_net_1 , 
        \un139_poly_mux[3]_net_1 , \un139_poly_mux[12]_net_1 , 
        \poly_mux_1[26]_net_1 , \un129_poly_mux[2]_net_1 , 
        \un129_poly_mux[1]_net_1 , \un129_poly_mux[10]_net_1 , 
        \crc_init_justified_1[31]_net_1 , 
        \crc_init_justified_0[31]_net_1 , \un1_crc_init_justified[6] , 
        \crc_init_justified_1[25]_net_1 , 
        \un30_crc_init_justified[1]_net_1 , 
        \un30_crc_init_justified[0]_net_1 , 
        \un30_crc_init_justified[9]_net_1 , 
        \crc_init_justified_1[30]_net_1 , 
        \un5_crc_init_justified[6]_net_1 , 
        \un5_crc_init_justified[5]_net_1 , 
        \un5_crc_init_justified[14]_net_1 , 
        \crc_init_justified_1[26]_net_1 , 
        \un25_crc_init_justified[2]_net_1 , 
        \un25_crc_init_justified[1]_net_1 , 
        \un25_crc_init_justified[10]_net_1 , 
        \crc_init_justified_1[29]_net_1 , 
        \crc_init_justified_0[29]_net_1 , 
        \un10_crc_init_justified[4]_net_1 , 
        \crc_init_justified[31]_net_1 , \poly_mux[26]_net_1 , 
        \un129_poly_mux[26]_net_1 , \poly_mux[25]_net_1 , 
        \un124_poly_mux[25]_net_1 , \poly_mux[30]_net_1 , 
        \poly_mux[29]_net_1 , \un144_poly_mux[13]_net_1 , 
        \un144_poly_mux[29]_net_1 , \un10_crc_out[26]_net_1 , 
        \un10_crc_out[27]_net_1 , \poly_mux[24]_net_1 , 
        \un119_poly_mux[8]_net_1 , \un119_poly_mux[0]_net_1 , 
        \un119_poly_mux[24]_net_1 , \crc_init_justified[24]_net_1 , 
        \un35_crc_init_justified[8]_net_1 , 
        \un35_crc_init_justified[0]_net_1 , 
        \un35_crc_init_justified[24]_net_1 , \crc_comb_out[8][31] , 
        \crc_comb_out[8][30] , \un30_crc_out[31]_net_1 , 
        \un30_crc_out[30]_net_1 , \poly_mux[28]_net_1 , 
        \un139_poly_mux[28]_net_1 , \un1_crc_out[16] , 
        \un1_crc_out[25] , \poly_mux[31]_net_1 , \un154_poly_mux[15] , 
        \un154_poly_mux[31] , \poly_mux[27]_net_1 , 
        \un134_poly_mux[11]_net_1 , \un134_poly_mux[27]_net_1 , 
        \un79_poly_mux[0]_net_1 , \un79_poly_mux[16]_net_1 , 
        \un84_poly_mux[1]_net_1 , \un84_poly_mux[17]_net_1 , 
        \un89_poly_mux[2]_net_1 , \un89_poly_mux[18]_net_1 , 
        \un130_crc_init_justified[5]_net_1 , 
        \un115_crc_init_justified[8]_net_1 , 
        \un105_crc_init_justified[10]_net_1 , 
        \un100_crc_init_justified[11]_net_1 , 
        \un95_crc_init_justified[12]_net_1 , 
        \un90_crc_init_justified[13]_net_1 , 
        \un85_crc_init_justified[14]_net_1 , 
        \un80_crc_init_justified[15]_net_1 , 
        \un75_crc_init_justified[0]_net_1 , 
        \un75_crc_init_justified[16]_net_1 , 
        \un70_crc_init_justified[1]_net_1 , 
        \un70_crc_init_justified[17]_net_1 , 
        \un65_crc_init_justified[2]_net_1 , 
        \un65_crc_init_justified[18]_net_1 , 
        \un60_crc_init_justified[3]_net_1 , 
        \un60_crc_init_justified[19]_net_1 , 
        \un50_crc_init_justified[21]_net_1 , 
        \un45_crc_init_justified[22]_net_1 , 
        \un30_crc_init_justified[25]_net_1 , 
        \un25_crc_init_justified[26]_net_1 , 
        \un20_crc_init_justified[27]_net_1 , 
        \un15_crc_init_justified[28]_net_1 , 
        \un10_crc_init_justified[29]_net_1 , 
        \crc_init_justified[22]_net_1 , \crc_init_justified[21]_net_1 , 
        \feedback[25] , \crc_in_masked[24] , \un45_crc_out[25]_net_1 , 
        \feedback[16] , \crc_in_masked[15] , \un109_poly_mux[6]_net_1 , 
        \un109_poly_mux[22]_net_1 , \feedback[21] , \crc_out_1_4[21] , 
        \feedback[22] , \crc_out_1_6[22] , \poly_mux[15] , 
        \un94_poly_mux[3]_net_1 , \un94_poly_mux[19]_net_1 , 
        \un99_poly_mux[4]_net_1 , \un99_poly_mux[20]_net_1 , 
        \un114_poly_mux[7]_net_1 , \un114_poly_mux[23]_net_1 , 
        \poly_mux[23]_net_1 , \poly_mux[13] , \crc_comb_out[8][19] , 
        \un15_crc_out[27]_net_1 , \crc_comb_out[8][27] , 
        \feedback[18] , \crc_out_1_1[18] , \un50_crc_out[10]_net_1 , 
        \feedback[10] , \crc_out_1_6[10] , \crc_comb_out[8][7] , 
        \poly_mux[12] , \crc_comb_out[8][13] , 
        \un65_crc_out[29]_net_1 , \un110_crc_init_justified[9]_net_1 , 
        \poly_mux[8] , \poly_mux[1] , \poly_mux[6] , 
        \un40_crc_out[8]_net_1 , \feedback[8] , \crc_out_1_6[8] , 
        \crc_comb_out[8][24] , \feedback[24] , 
        \crc_init_justified[23]_net_1 , 
        \un40_crc_init_justified[23]_net_1 , \poly_mux[10] , 
        \un70_crc_out[30]_net_1 , \crc_comb_out[8][14] , 
        \un5_crc_init_justified[30]_net_1 , \poly_mux[9] , 
        \un55_crc_out[11]_net_1 , \feedback[11] , \crc_out_1_6[11] , 
        \feedback[20] , \crc_out_1_3[20] , \un20_crc_out[20]_net_1 , 
        \un20_crc_out[4]_net_1 , \feedback[4] , \crc_out_1_2[4] , 
        \un104_poly_mux[21]_net_1 , \un104_poly_mux[5]_net_1 , 
        \un55_crc_init_justified[20]_net_1 , 
        \un55_crc_init_justified[4]_net_1 , \crc_comb_out[1][0] , 
        \feedback[13] , \feedback[14] , \feedback_0[25] , 
        \feedback_0[16] , \feedback[17] , \feedback_0[24] , 
        \feedback[3] , \feedback_0[18] , \feedback[19] , 
        \feedback_0[22] , \feedback_0[11] , \feedback_0[20] , 
        \feedback[2] , \feedback[7] , \feedback[31] , \feedback[5] , 
        \feedback[9] , \feedback_0[21] , N_170_0_0, N_170, 
        \crc_out_1_0[24] , \crc_in_masked_0[24] , 
        \crc_comb_out[2][23] , \crc_comb_out[2][15] , 
        \crc_comb_out[2][0] , \feedback_1[16] , \feedback_0[17] , 
        \feedback_1[18] , \feedback_0[19] , \feedback_1[20] , 
        \feedback_1[11] , \feedback[12] , \feedback_0[13] , 
        \feedback_0[7] , \feedback_0[10] , \feedback_0[4] , 
        \feedback_0[3] , \feedback_0[2] , \feedback_0[8] , 
        \feedback[6] , \feedback_1[21] , \feedback_0[5] , 
        \feedback_0[31] , \feedback_1[24] , \feedback_0[14] , 
        \feedback_1[22] , N_170_0_1, N_170_1, \crc_out_1_1[15] , 
        \crc_comb_out[3][23] , \crc_comb_out[3][24] , 
        \crc_in_masked_1[24] , \feedback_1[31] , \feedback_2[21] , 
        \feedback_1[13] , \feedback_1[14] , \feedback_2[22] , 
        \feedback_2[16] , \feedback_1[17] , \feedback_2[18] , 
        \feedback_1[19] , \feedback_2[20] , \feedback_2[11] , 
        \feedback_0[12] , \feedback[15] , \feedback_1[8] , 
        \feedback_1[5] , \feedback_1[2] , \feedback_1[4] , 
        \feedback_1[3] , \feedback_0[9] , \feedback_1[10] , 
        \feedback_1[7] , \feedback_0[6] , N_170_0_2, N_170_2, 
        \crc_out_1_2[23] , \crc_in_masked_0[15] , \feedback_2[31] , 
        \feedback_3[21] , \feedback_3[22] , \feedback_3[20] , 
        \feedback_2[13] , \feedback_2[14] , \feedback_1[25] , 
        \feedback_3[16] , \feedback_2[17] , \feedback_3[18] , 
        \feedback_2[19] , \feedback_1[12] , \feedback_1[6] , 
        \feedback_2[3] , \feedback[1] , \feedback_2[5] , 
        \feedback_2[4] , \feedback_2[10] , \feedback_3[11] , 
        \feedback_2[8] , \feedback[23] , \feedback_2[7] , 
        \crc_comb_out[4][15] , \crc_comb_out[4][24] , 
        \crc_comb_out[4][0] , N_170_0_3, N_170_3, \crc_out_1_3[15] , 
        \crc_in_masked[23] , \crc_in_masked_2[24] , 
        \crc_comb_out[5][23] , \crc_comb_out[5][0] , \feedback_3[31] , 
        \feedback_4[21] , \feedback_4[22] , \feedback_3[19] , 
        \feedback_4[20] , \feedback_3[13] , \feedback_3[14] , 
        \feedback_4[11] , \feedback_2[12] , \feedback_2[25] , 
        \feedback[26] , \feedback[28] , \feedback_2[24] , 
        \feedback_3[17] , \feedback_4[18] , \feedback_0[15] , 
        \feedback_3[7] , \feedback_3[4] , \feedback_2[2] , 
        \feedback_3[3] , \feedback_2[6] , \feedback_3[5] , 
        \feedback_1[9] , \feedback_4[16] , \feedback_3[8] , N_170_0_4, 
        N_170_4, \crc_out_1_4[23] , \crc_out_1_4[15] , 
        \crc_in_masked_1[15] , \crc_in_masked_3[24] , 
        \crc_comb_out[6][0] , \crc_comb_out[6][24] , \feedback_4[31] , 
        \feedback_5[21] , \feedback_5[18] , \feedback_4[19] , 
        \feedback_5[20] , \feedback_4[14] , \feedback_5[11] , 
        \feedback_5[22] , \feedback_3[12] , \feedback_1[15] , 
        \feedback_4[13] , \feedback[27] , \feedback[29] , 
        \feedback_0[23] , \feedback_3[25] , \feedback_5[16] , 
        \feedback_4[7] , \feedback_4[8] , \feedback_4[5] , 
        \feedback_4[3] , \feedback_4[4] , \feedback_3[6] , 
        \feedback_3[10] , \feedback_4[17] , \feedback_2[9] , 
        \feedback_3[2] , N_170_0_5, N_170_5, \crc_out_1_5[15] , 
        \crc_comb_out[7][0] , \crc_comb_out[7][23] , 
        \crc_in_masked_0[23] , \crc_in_masked_2[15] , \feedback_5[31] , 
        \feedback_6[21] , \feedback_6[22] , \feedback_5[17] , 
        \feedback_5[19] , \feedback_6[20] , \feedback_5[14] , 
        \feedback_3[9] , \feedback_4[12] , \feedback_5[13] , 
        \feedback_6[11] , \feedback_6[18] , \feedback_4[10] , 
        \feedback_0[26] , \feedback_0[28] , \feedback[30] , 
        \feedback_3[24] , \feedback_4[25] , \feedback_2[15] , 
        \feedback_5[8] , \feedback_0[1] , \feedback_4[6] , 
        \feedback_5[4] , \feedback_5[5] , \feedback_5[7] , 
        \feedback_6[16] , \feedback_4[2] , \feedback_5[3] , N_170_0_6, 
        GND, VCC;
    
    NOR2B \un25_crc_init_justified[1]  (.A(crc_init_mux[1]), .B(
        crc_poly_size_74), .Y(\un25_crc_init_justified[1]_net_1 ));
    NOR2B \un135_crc_out[27]  (.A(\crc_comb_out[8][27] ), .B(
        crc_poly_size_77), .Y(crc_unit_out[27]));
    OR3 \crc_init_justified_1[30]  (.A(
        \un5_crc_init_justified[6]_net_1 ), .B(
        \un5_crc_init_justified[5]_net_1 ), .C(
        \un5_crc_init_justified[14]_net_1 ), .Y(
        \crc_init_justified_1[30]_net_1 ));
    AND2 \un5_crc_out[26]  (.A(crc_poly_size_74), .B(
        \crc_comb_out[8][26] ), .Y(\un5_crc_out[26]_net_1 ));
    OR3 \poly_mux[27]  (.A(\poly_mux_0[27]_net_1 ), .B(
        \un134_poly_mux[11]_net_1 ), .C(\un134_poly_mux[27]_net_1 ), 
        .Y(\poly_mux[27]_net_1 ));
    NOR2B \un20_crc_init_justified[27]  (.A(crc_init_mux[27]), .B(
        crc_poly_size_77), .Y(\un20_crc_init_justified[27]_net_1 ));
    NOR2B \un139_poly_mux[3]  (.A(crc_poly_out[3]), .B(
        crc_poly_size_74), .Y(\un139_poly_mux[3]_net_1 ));
    NOR2B \genblk2[0].un1_crc_out[24]  (.A(\feedback[24] ), .B(
        crc_poly_size_75_0), .Y(\un1_crc_out[24] ));
    NOR2B \un155_crc_out[31]  (.A(\crc_comb_out[8][31] ), .B(
        crc_poly_size_77), .Y(crc_unit_out[31]));
    NOR2B \un119_poly_mux[8]  (.A(crc_poly_out[8]), .B(
        crc_poly_size_76), .Y(\un119_poly_mux[8]_net_1 ));
    \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_0  
        \genblk4[1].CRC_COMB  (.crc_out_1_0({\crc_out_1_0[24] }), 
        .un5_crc_init_justified({\un5_crc_init_justified[30]_net_1 }), 
        .crc_init_justified_1({\crc_init_justified_1[30]_net_1 }), 
        .crc_data_in({crc_data_in[6]}), .un90_crc_init_justified({
        \un90_crc_init_justified[13]_net_1 }), .crc_in_masked({
        \crc_in_masked_0[24] }), .crc_init_justified({
        \crc_init_justified[23]_net_1 , \crc_init_justified[22]_net_1 , 
        \crc_init_justified[21]_net_1 }), .un79_poly_mux_16(
        \un79_poly_mux[16]_net_1 ), .un79_poly_mux_0(
        \un79_poly_mux[0]_net_1 ), .un84_poly_mux_16(
        \un84_poly_mux[17]_net_1 ), .un84_poly_mux_0(
        \un84_poly_mux[1]_net_1 ), .un89_poly_mux_16(
        \un89_poly_mux[18]_net_1 ), .un89_poly_mux_0(
        \un89_poly_mux[2]_net_1 ), .un94_poly_mux_16(
        \un94_poly_mux[19]_net_1 ), .un94_poly_mux_0(
        \un94_poly_mux[3]_net_1 ), .un99_poly_mux_16(
        \un99_poly_mux[20]_net_1 ), .un99_poly_mux_0(
        \un99_poly_mux[4]_net_1 ), .\crc_comb_out[2]_23 (
        \crc_comb_out[2][23] ), .\crc_comb_out[2]_15 (
        \crc_comb_out[2][15] ), .\crc_comb_out[2]_0 (
        \crc_comb_out[2][0] ), .poly_mux_17(\poly_mux[23]_net_1 ), 
        .poly_mux_25(\poly_mux[31]_net_1 ), .poly_mux_18(
        \poly_mux[24]_net_1 ), .poly_mux_6(\poly_mux[12] ), 
        .poly_mux_7(\poly_mux[13] ), .poly_mux_9(\poly_mux[15] ), 
        .poly_mux_4(\poly_mux[10] ), .poly_mux_2(\poly_mux[8] ), 
        .poly_mux_0(\poly_mux[6] ), .un104_poly_mux_16(
        \un104_poly_mux[21]_net_1 ), .un104_poly_mux_0(
        \un104_poly_mux[5]_net_1 ), .feedback_29(\feedback[31] ), 
        .feedback_20(\feedback_0[22] ), .feedback_12(\feedback[14] ), 
        .feedback_22(\feedback_0[24] ), .feedback_14(\feedback_1[16] ), 
        .feedback_15(\feedback_0[17] ), .feedback_16(\feedback_1[18] ), 
        .feedback_17(\feedback_0[19] ), .feedback_18(\feedback_1[20] ), 
        .feedback_9(\feedback_1[11] ), .feedback_10(\feedback[12] ), 
        .feedback_11(\feedback_0[13] ), .feedback_5(\feedback_0[7] ), 
        .feedback_8(\feedback_0[10] ), .feedback_2(\feedback_0[4] ), 
        .feedback_1(\feedback_0[3] ), .feedback_0_d0(\feedback_0[2] ), 
        .feedback_6(\feedback_0[8] ), .feedback_4(\feedback[6] ), 
        .feedback_19(\feedback_1[21] ), .feedback_3(\feedback_0[5] ), 
        .crc_poly_out_11(crc_poly_out[11]), .crc_poly_out_14(
        crc_poly_out[14]), .crc_poly_out_7(crc_poly_out[7]), 
        .crc_poly_out_4(crc_poly_out[4]), .crc_poly_out_0(
        crc_poly_out[0]), .crc_poly_out_3(crc_poly_out[3]), 
        .crc_poly_out_2(crc_poly_out[2]), .crc_poly_out_5(
        crc_poly_out[5]), .feedback_0_17(\feedback_0[31] ), 
        .feedback_0_10(\feedback_1[24] ), .feedback_0_0(
        \feedback_0[14] ), .feedback_0_8(\feedback_1[22] ), 
        .un109_poly_mux_16(\un109_poly_mux[22]_net_1 ), 
        .un109_poly_mux_0(\un109_poly_mux[6]_net_1 ), .N_170_0(
        N_170_0_1), .N_170(N_170), .N_170_1(N_170_1), 
        .crc_poly_size_74_0(crc_poly_size_74_0), .crc_poly_size_77(
        crc_poly_size_77));
    NOR2B \un10_crc_out[27]  (.A(\crc_comb_out[8][27] ), .B(
        crc_poly_size_74), .Y(\un10_crc_out[27]_net_1 ));
    NOR2B \un119_poly_mux[0]  (.A(crc_poly_out[0]), .B(
        crc_poly_size_75), .Y(\un119_poly_mux[0]_net_1 ));
    NOR2B \un120_crc_out[24]  (.A(\crc_comb_out[8][24] ), .B(
        crc_poly_size_77), .Y(crc_unit_out[24]));
    AO1 \crc_out_1_0[0]  (.A(\un1_crc_out_0[0] ), .B(N_170_0), .C(
        \un1_crc_out[24] ), .Y(\crc_out_1_0[0]_net_1 ));
    AO1 \crc_out_1[10]  (.A(\crc_comb_out[8][26] ), .B(
        crc_poly_size_76_0), .C(\un50_crc_out[10]_net_1 ), .Y(
        crc_unit_out[10]));
    AO1 \poly_mux[30]  (.A(crc_poly_out[30]), .B(crc_poly_size_77), .C(
        \poly_mux_1[30]_net_1 ), .Y(\poly_mux[30]_net_1 ));
    NOR2B \genblk1[31].un154_poly_mux[15]  (.A(crc_poly_out[15]), .B(
        crc_poly_size_76_1), .Y(\un154_poly_mux[15] ));
    XA1 \crc_out_1_1_RNO[1]  (.A(\feedback[25] ), .B(
        \crc_in_masked[24] ), .C(crc_poly_size_75_0), .Y(
        \un5_crc_out[25] ));
    NOR2B \un104_poly_mux[5]  (.A(crc_poly_out[5]), .B(
        crc_poly_size_76_1), .Y(\un104_poly_mux[5]_net_1 ));
    XA1 \un20_crc_out[20]  (.A(\feedback[20] ), .B(\crc_out_1_3[20] ), 
        .C(crc_poly_size_76_0), .Y(\un20_crc_out[20]_net_1 ));
    AO1 \crc_out_1_1_RNO_0[1]  (.A(\crc_comb_out[8][17] ), .B(
        crc_poly_size_76_0), .C(\un5_crc_out[1]_net_1 ), .Y(
        \crc_out_1_0[1] ));
    XA1 \un40_crc_out[8]  (.A(\feedback[8] ), .B(\crc_out_1_6[8] ), .C(
        crc_poly_size_77), .Y(\un40_crc_out[8]_net_1 ));
    NOR2B \un94_poly_mux[19]  (.A(crc_poly_out[19]), .B(
        crc_poly_size_77), .Y(\un94_poly_mux[19]_net_1 ));
    XA1 \un90_crc_out[18]  (.A(\feedback[18] ), .B(\crc_out_1_1[18] ), 
        .C(crc_poly_size_77), .Y(crc_unit_out[18]));
    NOR2B \genblk1[31].un154_poly_mux[6]  (.A(crc_poly_out[6]), .B(
        crc_poly_size_74_0), .Y(\un154_poly_mux[6] ));
    NOR2B \un65_crc_init_justified[18]  (.A(crc_init_mux[18]), .B(
        crc_poly_size_77), .Y(\un65_crc_init_justified[18]_net_1 ));
    AO1 \crc_init_justified_0[31]  (.A(crc_init_mux[7]), .B(
        crc_poly_size_75_0), .C(\un1_crc_init_justified[6] ), .Y(
        \crc_init_justified_0[31]_net_1 ));
    NOR2B \un144_poly_mux[5]  (.A(crc_poly_out[5]), .B(
        crc_poly_size_75), .Y(\un144_poly_mux[5]_net_1 ));
    NOR2B \genblk2[0].un1_crc_out_0[0]  (.A(crc_poly_out[0]), .B(
        crc_poly_size_77), .Y(\un1_crc_out_0[0] ));
    NOR2B \un139_poly_mux[28]  (.A(crc_poly_out[28]), .B(
        crc_poly_size_77), .Y(\un139_poly_mux[28]_net_1 ));
    XA1 \un20_crc_out[4]  (.A(\feedback[4] ), .B(\crc_out_1_2[4] ), .C(
        crc_poly_size_77), .Y(\un20_crc_out[4]_net_1 ));
    NOR2B \un149_poly_mux[6]  (.A(crc_poly_out[6]), .B(
        crc_poly_size_75), .Y(\un149_poly_mux[6]_net_1 ));
    \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_4  
        \genblk4[5].CRC_COMB  (.un70_crc_init_justified_16(
        \un70_crc_init_justified[17]_net_1 ), 
        .un70_crc_init_justified_0(\un70_crc_init_justified[1]_net_1 ), 
        .crc_out_1_4_8(\crc_out_1_4[23] ), .crc_out_1_4_0(
        \crc_out_1_4[15] ), .un110_crc_init_justified({
        \un110_crc_init_justified[9]_net_1 }), 
        .un25_crc_init_justified({\un25_crc_init_justified[26]_net_1 })
        , .crc_init_justified_1({\crc_init_justified_1[26]_net_1 }), 
        .crc_data_in({crc_data_in[2]}), .crc_out_1_3({
        \crc_out_1_3[15] }), .crc_in_masked_0(\crc_in_masked_1[15] ), 
        .crc_in_masked_9(\crc_in_masked_3[24] ), .crc_in_masked_8(
        \crc_in_masked[23] ), .un104_poly_mux_16(
        \un104_poly_mux[21]_net_1 ), .un104_poly_mux_0(
        \un104_poly_mux[5]_net_1 ), .\crc_comb_out[6]_0 (
        \crc_comb_out[6][0] ), .\crc_comb_out[6]_24 (
        \crc_comb_out[6][24] ), .\crc_comb_out[5] ({
        \crc_comb_out[5][23] }), .un79_poly_mux_16(
        \un79_poly_mux[16]_net_1 ), .un79_poly_mux_0(
        \un79_poly_mux[0]_net_1 ), .un89_poly_mux_16(
        \un89_poly_mux[18]_net_1 ), .un89_poly_mux_0(
        \un89_poly_mux[2]_net_1 ), .un94_poly_mux_16(
        \un94_poly_mux[19]_net_1 ), .un94_poly_mux_0(
        \un94_poly_mux[3]_net_1 ), .un99_poly_mux_16(
        \un99_poly_mux[20]_net_1 ), .un99_poly_mux_0(
        \un99_poly_mux[4]_net_1 ), .un109_poly_mux_16(
        \un109_poly_mux[22]_net_1 ), .un109_poly_mux_0(
        \un109_poly_mux[6]_net_1 ), .feedback_0_20(\feedback_4[31] ), 
        .feedback_0_10(\feedback_5[21] ), .feedback_0_7(
        \feedback_5[18] ), .feedback_0_8(\feedback_4[19] ), 
        .feedback_0_9(\feedback_5[20] ), .feedback_0_3(
        \feedback_4[14] ), .feedback_0_0(\feedback_5[11] ), 
        .feedback_0_11(\feedback_5[22] ), .feedback_0_1(
        \feedback_3[12] ), .feedback_0_4(\feedback_1[15] ), 
        .feedback_0_2(\feedback_4[13] ), .un84_poly_mux_16(
        \un84_poly_mux[17]_net_1 ), .un84_poly_mux_0(
        \un84_poly_mux[1]_net_1 ), .poly_mux_4(\poly_mux[10] ), 
        .poly_mux_24(\poly_mux[30]_net_1 ), .poly_mux_23(
        \poly_mux[29]_net_1 ), .poly_mux_22(\poly_mux[28]_net_1 ), 
        .poly_mux_21(\poly_mux[27]_net_1 ), .poly_mux_25(
        \poly_mux[31]_net_1 ), .poly_mux_17(\poly_mux[23]_net_1 ), 
        .poly_mux_18(\poly_mux[24]_net_1 ), .poly_mux_19(
        \poly_mux[25]_net_1 ), .poly_mux_2(\poly_mux[8] ), .poly_mux_0(
        \poly_mux[6] ), .poly_mux_9(\poly_mux[15] ), .poly_mux_7(
        \poly_mux[13] ), .poly_mux_3(\poly_mux[9] ), .feedback_29(
        \feedback_3[31] ), .feedback_19(\feedback_3[21] ), 
        .feedback_20(\feedback_4[22] ), .feedback_17(\feedback_0[19] ), 
        .feedback_18(\feedback_2[20] ), .feedback_16(\feedback_0[18] ), 
        .feedback_11(\feedback_2[13] ), .feedback_12(\feedback_3[14] ), 
        .feedback_9(\feedback_1[11] ), .feedback_10(\feedback_0[12] ), 
        .feedback_13(\feedback_0[15] ), .feedback_22(\feedback_2[24] ), 
        .feedback_25(\feedback[27] ), .feedback_27(\feedback[29] ), 
        .feedback_21(\feedback_0[23] ), .feedback_23(\feedback_3[25] ), 
        .feedback_14(\feedback_5[16] ), .feedback_5(\feedback_4[7] ), 
        .feedback_6(\feedback_4[8] ), .feedback_3(\feedback_4[5] ), 
        .feedback_1(\feedback_4[3] ), .feedback_2(\feedback_4[4] ), 
        .feedback_4(\feedback_3[6] ), .feedback_8(\feedback_3[10] ), 
        .feedback_15(\feedback_4[17] ), .feedback_7(\feedback_2[9] ), 
        .feedback_0_d0(\feedback_3[2] ), .crc_poly_out_0(
        crc_poly_out[0]), .crc_poly_out_14(crc_poly_out[14]), 
        .crc_poly_out_7(crc_poly_out[7]), .crc_poly_out_5(
        crc_poly_out[5]), .crc_poly_out_11(crc_poly_out[11]), 
        .crc_poly_out_3(crc_poly_out[3]), .crc_poly_out_4(
        crc_poly_out[4]), .crc_poly_out_12(crc_poly_out[12]), 
        .crc_poly_out_10(crc_poly_out[10]), .crc_poly_out_2(
        crc_poly_out[2]), .N_170_0(N_170_0_5), .N_170_0_0(N_170_0_0), 
        .N_170_0_1(N_170_0_3), .N_170(N_170_2), .N_170_0_2(N_170_0_1), 
        .N_170_1(N_170_5), .crc_poly_size_76_1(crc_poly_size_76_1), 
        .crc_poly_size_74_0(crc_poly_size_74_0), .crc_poly_size_75_0(
        crc_poly_size_75_0), .crc_poly_size_77(crc_poly_size_77));
    AO1 \crc_out_1_0[5]  (.A(\crc_comb_out[8][5] ), .B(
        crc_poly_size_77), .C(\un25_crc_out[21]_net_1 ), .Y(
        \crc_out_1_0[5]_net_1 ));
    NOR2B \un139_poly_mux[12]  (.A(crc_poly_out[12]), .B(
        crc_poly_size_76), .Y(\un139_poly_mux[12]_net_1 ));
    NOR2B \un114_poly_mux[7]  (.A(crc_poly_out[7]), .B(
        crc_poly_size_76_1), .Y(\un114_poly_mux[7]_net_1 ));
    NOR2B \un5_crc_init_justified[30]  (.A(crc_init_mux[30]), .B(
        crc_poly_size_77), .Y(\un5_crc_init_justified[30]_net_1 ));
    NOR2B \un40_crc_init_justified[23]  (.A(crc_init_mux[23]), .B(
        crc_poly_size_77), .Y(\un40_crc_init_justified[23]_net_1 ));
    NOR2B \un84_poly_mux[17]  (.A(crc_poly_out[17]), .B(
        crc_poly_size_77), .Y(\un84_poly_mux[17]_net_1 ));
    NOR2B \un15_crc_out[27]  (.A(\crc_comb_out[8][27] ), .B(
        crc_poly_size_75), .Y(\un15_crc_out[27]_net_1 ));
    NOR2B \un39_poly_mux[8]  (.A(crc_poly_out[8]), .B(crc_poly_size_77)
        , .Y(\poly_mux[8] ));
    NOR2B \crc_init_justified_0_RNO_0[27]  (.A(crc_init_mux[2]), .B(
        crc_poly_size_74_0), .Y(\un20_crc_init_justified[2] ));
    OR3 \poly_mux_1[26]  (.A(\un129_poly_mux[2]_net_1 ), .B(
        \un129_poly_mux[1]_net_1 ), .C(\un129_poly_mux[10]_net_1 ), .Y(
        \poly_mux_1[26]_net_1 ));
    OR2 \crc_init_justified_0[28]  (.A(\un15_crc_init_justified[4] ), 
        .B(\un15_crc_init_justified[3] ), .Y(
        \crc_init_justified_0[28]_net_1 ));
    NOR2B \un30_crc_init_justified[0]  (.A(crc_init_mux[0]), .B(
        crc_poly_size_74), .Y(\un30_crc_init_justified[0]_net_1 ));
    NOR2B \un115_crc_out[23]  (.A(\crc_comb_out[8][23] ), .B(
        crc_poly_size_77), .Y(crc_unit_out[23]));
    OR3 \poly_mux[24]  (.A(\un119_poly_mux[8]_net_1 ), .B(
        \un119_poly_mux[0]_net_1 ), .C(\un119_poly_mux[24]_net_1 ), .Y(
        \poly_mux[24]_net_1 ));
    NOR2B \un30_crc_out[31]  (.A(\crc_comb_out[8][31] ), .B(
        crc_poly_size_74), .Y(\un30_crc_out[31]_net_1 ));
    AO1 \crc_init_justified[22]  (.A(crc_init_mux[6]), .B(
        crc_poly_size_76_0), .C(\un45_crc_init_justified[22]_net_1 ), 
        .Y(\crc_init_justified[22]_net_1 ));
    NOR2B \un104_poly_mux[21]  (.A(crc_poly_out[21]), .B(
        crc_poly_size_77), .Y(\un104_poly_mux[21]_net_1 ));
    GND GND_i (.Y(GND));
    OR2 \crc_init_justified_0[27]  (.A(\un20_crc_init_justified[3] ), 
        .B(\un20_crc_init_justified[2] ), .Y(
        \crc_init_justified_0[27]_net_1 ));
    NOR2B \un99_poly_mux[4]  (.A(crc_poly_out[4]), .B(crc_poly_size_76)
        , .Y(\un99_poly_mux[4]_net_1 ));
    NOR2B \un129_poly_mux[26]  (.A(crc_poly_out[26]), .B(
        crc_poly_size_77), .Y(\un129_poly_mux[26]_net_1 ));
    AO1 \crc_out_1[11]  (.A(\crc_comb_out[8][27] ), .B(
        crc_poly_size_76_0), .C(\un55_crc_out[11]_net_1 ), .Y(
        crc_unit_out[11]));
    NOR2B \un139_poly_mux[4]  (.A(crc_poly_out[4]), .B(
        crc_poly_size_75), .Y(\un139_poly_mux[4]_net_1 ));
    XA1 \un110_crc_out[22]  (.A(\feedback[22] ), .B(\crc_out_1_6[22] ), 
        .C(crc_poly_size_77), .Y(crc_unit_out[22]));
    OR3 \poly_mux_1[25]  (.A(\un124_poly_mux[1]_net_1 ), .B(
        \un124_poly_mux[0]_net_1 ), .C(\un124_poly_mux[9]_net_1 ), .Y(
        \poly_mux_1[25]_net_1 ));
    \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_3  
        \genblk4[4].CRC_COMB  (.\crc_comb_out[4] ({
        \crc_comb_out[4][24] }), .crc_out_1_3({\crc_out_1_3[15] }), 
        .un105_crc_init_justified({
        \un105_crc_init_justified[10]_net_1 }), 
        .un65_crc_init_justified_16(
        \un65_crc_init_justified[18]_net_1 ), 
        .un65_crc_init_justified_0(\un65_crc_init_justified[2]_net_1 ), 
        .un20_crc_init_justified({\un20_crc_init_justified[27]_net_1 })
        , .crc_init_justified_1({\crc_init_justified_1[27]_net_1 }), 
        .crc_data_in({crc_data_in[3]}), .crc_in_masked({
        \crc_in_masked_2[24] , \crc_in_masked[23] }), .crc_out_1_2_0({
        \crc_out_1_2[23] }), .\crc_comb_out[5]_23 (
        \crc_comb_out[5][23] ), .\crc_comb_out[5]_0 (
        \crc_comb_out[5][0] ), .un104_poly_mux_16(
        \un104_poly_mux[21]_net_1 ), .un104_poly_mux_0(
        \un104_poly_mux[5]_net_1 ), .un109_poly_mux_16(
        \un109_poly_mux[22]_net_1 ), .un109_poly_mux_0(
        \un109_poly_mux[6]_net_1 ), .un84_poly_mux_16(
        \un84_poly_mux[17]_net_1 ), .un84_poly_mux_0(
        \un84_poly_mux[1]_net_1 ), .un89_poly_mux_16(
        \un89_poly_mux[18]_net_1 ), .un89_poly_mux_0(
        \un89_poly_mux[2]_net_1 ), .un94_poly_mux_16(
        \un94_poly_mux[19]_net_1 ), .un94_poly_mux_0(
        \un94_poly_mux[3]_net_1 ), .un99_poly_mux_16(
        \un99_poly_mux[20]_net_1 ), .un99_poly_mux_0(
        \un99_poly_mux[4]_net_1 ), .feedback_0_12(\feedback[23] ), 
        .feedback_0_20(\feedback_3[31] ), .feedback_0_10(
        \feedback_4[21] ), .feedback_0_11(\feedback_4[22] ), 
        .feedback_0_8(\feedback_3[19] ), .feedback_0_9(
        \feedback_4[20] ), .feedback_0_2(\feedback_3[13] ), 
        .feedback_0_3(\feedback_3[14] ), .feedback_0_0(
        \feedback_4[11] ), .feedback_0_1(\feedback_2[12] ), 
        .crc_poly_out_0(crc_poly_out[0]), .crc_poly_out_14(
        crc_poly_out[14]), .crc_poly_out_7(crc_poly_out[7]), 
        .crc_poly_out_4(crc_poly_out[4]), .crc_poly_out_2(
        crc_poly_out[2]), .crc_poly_out_3(crc_poly_out[3]), 
        .crc_poly_out_5(crc_poly_out[5]), .crc_poly_out_11(
        crc_poly_out[11]), .crc_poly_out_9(crc_poly_out[9]), 
        .un79_poly_mux_16(\un79_poly_mux[16]_net_1 ), .un79_poly_mux_0(
        \un79_poly_mux[0]_net_1 ), .feedback_29(\feedback_2[31] ), 
        .feedback_23(\feedback_2[25] ), .feedback_11(\feedback_1[13] ), 
        .feedback_12(\feedback_2[14] ), .feedback_9(\feedback_0[11] ), 
        .feedback_10(\feedback[12] ), .feedback_18(\feedback_1[20] ), 
        .feedback_19(\feedback_2[21] ), .feedback_17(\feedback[19] ), 
        .feedback_20(\feedback_3[22] ), .feedback_24(\feedback[26] ), 
        .feedback_26(\feedback[28] ), .feedback_22(\feedback_2[24] ), 
        .feedback_15(\feedback_3[17] ), .feedback_16(\feedback_4[18] ), 
        .feedback_13(\feedback_0[15] ), .feedback_5(\feedback_3[7] ), 
        .feedback_2(\feedback_3[4] ), .feedback_0_d0(\feedback_2[2] ), 
        .feedback_1(\feedback_3[3] ), .feedback_4(\feedback_2[6] ), 
        .feedback_3(\feedback_3[5] ), .feedback_7(\feedback_1[9] ), 
        .feedback_14(\feedback_4[16] ), .feedback_6(\feedback_3[8] ), 
        .poly_mux_19(\poly_mux[25]_net_1 ), .poly_mux_24(
        \poly_mux[30]_net_1 ), .poly_mux_23(\poly_mux[29]_net_1 ), 
        .poly_mux_22(\poly_mux[28]_net_1 ), .poly_mux_20(
        \poly_mux[26]_net_1 ), .poly_mux_25(\poly_mux[31]_net_1 ), 
        .poly_mux_17(\poly_mux[23]_net_1 ), .poly_mux_18(
        \poly_mux[24]_net_1 ), .poly_mux_7(\poly_mux[13] ), 
        .poly_mux_9(\poly_mux[15] ), .poly_mux_0(\poly_mux[6] ), 
        .poly_mux_6(\poly_mux[12] ), .poly_mux_2(\poly_mux[8] ), 
        .N_170_0(N_170_0_4), .crc_poly_size_74(crc_poly_size_74), 
        .N_170(N_170_4), .N_170_0_0(N_170_0_2), .N_170_0_1(N_170_0_1), 
        .N_170_0_2(N_170_0_0), .crc_poly_size_75_0(crc_poly_size_75_0), 
        .crc_poly_size_77(crc_poly_size_77));
    XA1 \un10_crc_out[18]  (.A(\feedback[18] ), .B(\crc_out_1_1[18] ), 
        .C(crc_poly_size_76_0), .Y(\un10_crc_out[18]_net_1 ));
    NOR2B \un79_poly_mux[16]  (.A(crc_poly_out[16]), .B(
        crc_poly_size_77), .Y(\un79_poly_mux[16]_net_1 ));
    AO1 \crc_init_justified_1[31]  (.A(crc_init_mux[15]), .B(
        crc_poly_size_76_0), .C(\crc_init_justified_0[31]_net_1 ), .Y(
        \crc_init_justified_1[31]_net_1 ));
    XA1 \un30_crc_out[22]  (.A(\feedback[22] ), .B(\crc_out_1_6[22] ), 
        .C(crc_poly_size_76_0), .Y(\un30_crc_out[22]_net_1 ));
    NOR2B \crc_init_justified_0_RNO_0[28]  (.A(crc_init_mux[3]), .B(
        crc_poly_size_74), .Y(\un15_crc_init_justified[3] ));
    XA1 \genblk2[0].un1_crc_out[25]  (.A(\feedback[25] ), .B(
        \crc_in_masked[24] ), .C(crc_poly_size_74_0), .Y(
        \un1_crc_out[25] ));
    NOR2B \un10_crc_out[26]  (.A(\crc_comb_out[8][26] ), .B(
        crc_poly_size_75), .Y(\un10_crc_out[26]_net_1 ));
    NOR2B \genblk1[31].un154_poly_mux[31]  (.A(crc_poly_out[31]), .B(
        crc_poly_size_77), .Y(\un154_poly_mux[31] ));
    NOR2B \un144_poly_mux[13]  (.A(crc_poly_out[13]), .B(
        crc_poly_size_76_1), .Y(\un144_poly_mux[13]_net_1 ));
    AO1 \crc_out_1[5]  (.A(\crc_comb_out[8][30] ), .B(
        crc_poly_size_74_0), .C(\crc_out_1_1[5]_net_1 ), .Y(
        crc_unit_out[5]));
    NOR2B \un5_crc_init_justified[14]  (.A(crc_init_mux[14]), .B(
        crc_poly_size_76), .Y(\un5_crc_init_justified[14]_net_1 ));
    NOR2B \un10_crc_init_justified[29]  (.A(crc_init_mux[29]), .B(
        crc_poly_size_77), .Y(\un10_crc_init_justified[29]_net_1 ));
    NOR2B \un84_poly_mux[1]  (.A(crc_poly_out[1]), .B(
        crc_poly_size_76_1), .Y(\un84_poly_mux[1]_net_1 ));
    AO1 \poly_mux_0[27]  (.A(crc_poly_out[2]), .B(crc_poly_size_74_0), 
        .C(\un134_poly_mux[3]_net_1 ), .Y(\poly_mux_0[27]_net_1 ));
    NOR2B \un75_crc_init_justified[0]  (.A(crc_init_mux[0]), .B(
        crc_poly_size_76_1), .Y(\un75_crc_init_justified[0]_net_1 ));
    NOR2B \un114_poly_mux[23]  (.A(crc_poly_out[23]), .B(
        crc_poly_size_77), .Y(\un114_poly_mux[23]_net_1 ));
    OR2 \crc_init_justified_1[28]  (.A(
        \crc_init_justified_0[28]_net_1 ), .B(
        \un15_crc_init_justified[12]_net_1 ), .Y(
        \crc_init_justified_1[28]_net_1 ));
    NOR2B \un130_crc_init_justified[5]  (.A(crc_init_mux[5]), .B(
        crc_poly_size_77), .Y(\un130_crc_init_justified[5]_net_1 ));
    NOR2B \un115_crc_init_justified[8]  (.A(crc_init_mux[8]), .B(
        crc_poly_size_77), .Y(\un115_crc_init_justified[8]_net_1 ));
    NOR2B \un85_crc_out[17]  (.A(\crc_comb_out[8][17] ), .B(
        crc_poly_size_77), .Y(crc_unit_out[17]));
    XA1 \un100_crc_out[20]  (.A(\feedback[20] ), .B(\crc_out_1_3[20] ), 
        .C(crc_poly_size_77), .Y(crc_unit_out[20]));
    NOR2B \un100_crc_init_justified[11]  (.A(crc_init_mux[11]), .B(
        crc_poly_size_77), .Y(\un100_crc_init_justified[11]_net_1 ));
    AO1 \poly_mux_0[29]  (.A(crc_poly_out[4]), .B(crc_poly_size_74_0), 
        .C(\un144_poly_mux[5]_net_1 ), .Y(\poly_mux_0[29]_net_1 ));
    OR2 \poly_mux[28]  (.A(\poly_mux_1[28]_net_1 ), .B(
        \un139_poly_mux[28]_net_1 ), .Y(\poly_mux[28]_net_1 ));
    OR2 \crc_init_justified_1[27]  (.A(
        \crc_init_justified_0[27]_net_1 ), .B(
        \un20_crc_init_justified[11]_net_1 ), .Y(
        \crc_init_justified_1[27]_net_1 ));
    OR2 \poly_mux[26]  (.A(\poly_mux_1[26]_net_1 ), .B(
        \un129_poly_mux[26]_net_1 ), .Y(\poly_mux[26]_net_1 ));
    NOR2B \un30_crc_out[30]  (.A(\crc_comb_out[8][30] ), .B(
        crc_poly_size_75), .Y(\un30_crc_out[30]_net_1 ));
    VCC VCC_i (.Y(VCC));
    NOR2B \un129_poly_mux[1]  (.A(crc_poly_out[1]), .B(
        crc_poly_size_74), .Y(\un129_poly_mux[1]_net_1 ));
    NOR2B \un134_poly_mux[3]  (.A(crc_poly_out[3]), .B(
        crc_poly_size_75), .Y(\un134_poly_mux[3]_net_1 ));
    OR3 \poly_mux_1[28]  (.A(\un139_poly_mux[4]_net_1 ), .B(
        \un139_poly_mux[3]_net_1 ), .C(\un139_poly_mux[12]_net_1 ), .Y(
        \poly_mux_1[28]_net_1 ));
    XA1 \un25_crc_out[21]  (.A(\feedback[21] ), .B(\crc_out_1_4[21] ), 
        .C(crc_poly_size_76_1), .Y(\un25_crc_out[21]_net_1 ));
    \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_6  
        \genblk4[7].CRC_COMB  (.un20_crc_out_16(
        \un20_crc_out[20]_net_1 ), .un20_crc_out_0(
        \un20_crc_out[4]_net_1 ), .\crc_comb_out[3] ({
        \crc_comb_out[3][24] }), .un85_crc_init_justified({
        \un85_crc_init_justified[14]_net_1 }), .crc_out_1_4_14(
        \crc_out_1_4[21] ), .un80_crc_init_justified({
        \un80_crc_init_justified[15]_net_1 }), .crc_out_1_3_14(
        \crc_out_1_3[20] ), .un130_crc_init_justified({
        \un130_crc_init_justified[5]_net_1 }), .\crc_comb_out[1] ({
        \crc_comb_out[1][0] }), .crc_out_1_6_14(\crc_out_1_6[22] ), 
        .crc_out_1_6_2(\crc_out_1_6[10] ), .crc_out_1_6_0(
        \crc_out_1_6[8] ), .crc_out_1_6_3(\crc_out_1_6[11] ), 
        .crc_out_1_2_0(\crc_out_1_2[4] ), .\crc_comb_out[4]_15 (
        \crc_comb_out[4][15] ), .\crc_comb_out[4]_0 (
        \crc_comb_out[4][0] ), .\crc_comb_out[2]_15 (
        \crc_comb_out[2][15] ), .\crc_comb_out[2]_0 (
        \crc_comb_out[2][0] ), .crc_out_1_1_14(\crc_out_1_1[18] ), 
        .crc_in_masked_0_9(\crc_in_masked_0[24] ), .crc_in_masked_0_0(
        \crc_in_masked_1[15] ), .\crc_comb_out[5] ({
        \crc_comb_out[5][0] }), .crc_init_justified({
        \crc_init_justified[24]_net_1 }), .crc_data_in({crc_data_in[0]})
        , .\crc_comb_out[6]_24 (\crc_comb_out[6][24] ), 
        .\crc_comb_out[6]_0 (\crc_comb_out[6][0] ), .un15_crc_out_0(
        \un15_crc_out[27]_net_1 ), .crc_out_1_0_0({
        \crc_out_1_0[3]_net_1 }), .crc_in_masked_1_9(
        \crc_in_masked_1[24] ), .crc_in_masked_1_0(
        \crc_in_masked_2[15] ), .crc_in_masked_2_9(
        \crc_in_masked_3[24] ), .crc_in_masked_2_0(\crc_in_masked[15] )
        , .crc_out_1_5_0({\crc_out_1_5[15] }), .crc_in_masked_3({
        \crc_in_masked[24] }), .feedback_30(\feedback_5[31] ), 
        .feedback_24(\feedback_2[25] ), .feedback_13(\feedback_5[14] ), 
        .feedback_12(\feedback_4[13] ), .feedback_11(\feedback_2[12] ), 
        .feedback_7(\feedback_5[8] ), .feedback_27(\feedback[28] ), 
        .feedback_28(\feedback[29] ), .feedback_25(\feedback[26] ), 
        .feedback_26(\feedback[27] ), .feedback_19(\feedback_5[20] ), 
        .feedback_20(\feedback_6[21] ), .feedback_17(\feedback_3[18] ), 
        .feedback_18(\feedback_3[19] ), .feedback_15(\feedback_1[16] ), 
        .feedback_16(\feedback_1[17] ), .feedback_10(\feedback_4[11] ), 
        .feedback_9(\feedback_2[10] ), .feedback_6_d0(\feedback[7] ), 
        .feedback_5_d0(\feedback_1[6] ), .feedback_3_d0(
        \feedback_0[4] ), .feedback_4_d0(\feedback_1[5] ), 
        .feedback_2_d0(\feedback[3] ), .feedback_1_d0(\feedback_2[2] ), 
        .feedback_21(\feedback_6[22] ), .feedback_23(\feedback_3[24] ), 
        .crc_in_masked_9(\crc_in_masked_2[24] ), .crc_in_masked_0_d0(
        \crc_in_masked_0[15] ), .crc_in_masked_8(\crc_in_masked_0[23] )
        , .feedback_1_24(\feedback_3[25] ), .feedback_1_16(
        \feedback_4[17] ), .feedback_1_17(\feedback_6[18] ), 
        .feedback_1_15(\feedback_4[16] ), .feedback_1_19(
        \feedback_4[20] ), .feedback_1_18(\feedback_2[19] ), 
        .feedback_1_7(\feedback_4[8] ), .feedback_1_8(\feedback_3[9] ), 
        .feedback_1_10(\feedback_5[11] ), .feedback_1_11(
        \feedback_4[12] ), .feedback_1_6(\feedback_0[7] ), 
        .feedback_1_2(\feedback_2[3] ), .feedback_1_3(\feedback_1[4] ), 
        .feedback_1_4(\feedback_2[5] ), .feedback_1_1(\feedback[2] ), 
        .feedback_1_9(\feedback_3[10] ), .feedback_1_5(\feedback[6] ), 
        .feedback_1_0(\feedback_0[1] ), .feedback_1_20(\feedback[21] ), 
        .un104_poly_mux_16(\un104_poly_mux[21]_net_1 ), 
        .un104_poly_mux_0(\un104_poly_mux[5]_net_1 ), 
        .un109_poly_mux_16(\un109_poly_mux[22]_net_1 ), 
        .un109_poly_mux_0(\un109_poly_mux[6]_net_1 ), .feedback_6_2(
        \feedback_5[5] ), .feedback_6_13(\feedback[16] ), 
        .un79_poly_mux_16(\un79_poly_mux[16]_net_1 ), .un79_poly_mux_0(
        \un79_poly_mux[0]_net_1 ), .feedback_4_5(\feedback_5[7] ), 
        .feedback_4_6(\feedback_3[8] ), .feedback_4_3(\feedback_0[5] ), 
        .feedback_4_1(\feedback_5[3] ), .feedback_4_14(
        \feedback_5[16] ), .feedback_4_15(\feedback_5[17] ), 
        .feedback_4_4(\feedback_4[6] ), .feedback_4_2(\feedback_5[4] ), 
        .feedback_4_23(\feedback[25] ), .feedback_4_16(\feedback[18] ), 
        .un89_poly_mux_16(\un89_poly_mux[18]_net_1 ), .un89_poly_mux_0(
        \un89_poly_mux[2]_net_1 ), .feedback_2_23(\feedback_4[25] ), 
        .feedback_2_16(\feedback_2[18] ), .feedback_2_14(
        \feedback_0[16] ), .feedback_2_15(\feedback_0[17] ), 
        .feedback_2_17(\feedback_5[19] ), .feedback_2_6(
        \feedback_1[8] ), .feedback_2_5(\feedback_4[7] ), 
        .feedback_2_1(\feedback_0[3] ), .feedback_2_7(\feedback_1[9] ), 
        .feedback_2_3(\feedback[5] ), .feedback_2_4(\feedback_3[6] ), 
        .feedback_2_2(\feedback_2[4] ), .feedback_2_0(\feedback_0[2] ), 
        .feedback_2_8(\feedback_4[10] ), .feedback_2_9(
        \feedback_6[11] ), .feedback_2_18(\feedback[20] ), 
        .un99_poly_mux_16(\un99_poly_mux[20]_net_1 ), .un99_poly_mux_0(
        \un99_poly_mux[4]_net_1 ), .un45_crc_out({
        \un45_crc_out[25]_net_1 }), .crc_init_mux_6(crc_init_mux[6]), 
        .crc_init_mux_2(crc_init_mux[2]), .crc_init_mux_4(
        crc_init_mux[4]), .crc_init_mux_0(crc_init_mux[0]), 
        .crc_init_mux_3(crc_init_mux[3]), .crc_init_mux_1(
        crc_init_mux[1]), .crc_init_mux_7(crc_init_mux[7]), 
        .\crc_comb_out[8]_0 (\crc_comb_out[8][1] ), 
        .\crc_comb_out[8]_14 (\crc_comb_out[8][15] ), 
        .\crc_comb_out[8]_25 (\crc_comb_out[8][26] ), 
        .\crc_comb_out[8]_26 (\crc_comb_out[8][27] ), 
        .\crc_comb_out[8]_28 (\crc_comb_out[8][29] ), 
        .\crc_comb_out[8]_29 (\crc_comb_out[8][30] ), 
        .\crc_comb_out[8]_30 (\crc_comb_out[8][31] ), 
        .\crc_comb_out[8]_22 (\crc_comb_out[8][23] ), 
        .\crc_comb_out[8]_1 (\crc_comb_out[8][2] ), 
        .\crc_comb_out[8]_6 (\crc_comb_out[8][7] ), 
        .\crc_comb_out[8]_12 (\crc_comb_out[8][13] ), 
        .\crc_comb_out[8]_4 (\crc_comb_out[8][5] ), 
        .\crc_comb_out[8]_5 (\crc_comb_out[8][6] ), 
        .\crc_comb_out[8]_13 (\crc_comb_out[8][14] ), 
        .\crc_comb_out[8]_16 (\crc_comb_out[8][17] ), 
        .\crc_comb_out[8]_2 (\crc_comb_out[8][3] ), 
        .\crc_comb_out[8]_18 (\crc_comb_out[8][19] ), 
        .\crc_comb_out[8]_23 (\crc_comb_out[8][24] ), 
        .\crc_comb_out[7]_0 (\crc_comb_out[7][0] ), 
        .\crc_comb_out[7]_23 (\crc_comb_out[7][23] ), .feedback_0_24(
        \feedback_1[25] ), .feedback_0_25(\feedback_0[26] ), 
        .feedback_0_18(\feedback_4[19] ), .feedback_0_19(
        \feedback_6[20] ), .feedback_0_16(\feedback_2[17] ), 
        .feedback_0_17(\feedback_4[18] ), .feedback_0_15(
        \feedback_2[16] ), .feedback_0_20(\feedback_5[21] ), 
        .feedback_0_11(\feedback_3[12] ), .feedback_0_8(
        \feedback_0[9] ), .feedback_0_7(\feedback_0[8] ), 
        .feedback_0_6(\feedback_3[7] ), .feedback_0_9(\feedback_1[10] )
        , .feedback_0_10(\feedback_3[11] ), .feedback_0_2(
        \feedback_4[3] ), .feedback_0_0(\feedback[1] ), .feedback_0_3(
        \feedback_3[4] ), .feedback_0_4(\feedback_4[5] ), 
        .feedback_0_1(\feedback_1[2] ), .feedback_0_5(\feedback_2[6] ), 
        .feedback_0_27(\feedback_0[28] ), .feedback_0_29(
        \feedback[30] ), .feedback_0_12(\feedback_5[13] ), 
        .feedback_0_14(\feedback_2[15] ), .feedback_0_21(
        \feedback[22] ), .feedback_0_23(\feedback[24] ), 
        .un84_poly_mux_16(\un84_poly_mux[17]_net_1 ), .un84_poly_mux_0(
        \un84_poly_mux[1]_net_1 ), .poly_mux_8(\poly_mux[9] ), 
        .poly_mux_26(\poly_mux[27]_net_1 ), .poly_mux_25(
        \poly_mux[26]_net_1 ), .poly_mux_24(\poly_mux[25]_net_1 ), 
        .poly_mux_28(\poly_mux[29]_net_1 ), .poly_mux_27(
        \poly_mux[28]_net_1 ), .poly_mux_14(\poly_mux[15] ), 
        .poly_mux_7(\poly_mux[8] ), .poly_mux_9(\poly_mux[10] ), 
        .poly_mux_5(\poly_mux[6] ), .poly_mux_0(\poly_mux[1] ), 
        .poly_mux_29(\poly_mux[30]_net_1 ), .poly_mux_12(
        \poly_mux[13] ), .poly_mux_30(\poly_mux[31]_net_1 ), 
        .poly_mux_22(\poly_mux[23]_net_1 ), .poly_mux_23(
        \poly_mux[24]_net_1 ), .poly_mux_11(\poly_mux[12] ), 
        .crc_unit_out_0(crc_unit_out[3]), .crc_unit_out_1(
        crc_unit_out[4]), .crc_unit_out_6(crc_unit_out[9]), 
        .crc_unit_out_25(crc_unit_out[28]), .crc_unit_out_9(
        crc_unit_out[12]), .un94_poly_mux_16(\un94_poly_mux[19]_net_1 )
        , .un94_poly_mux_0(\un94_poly_mux[3]_net_1 ), .feedback_3_16(
        \feedback_5[18] ), .feedback_3_14(\feedback_3[16] ), 
        .feedback_3_15(\feedback_3[17] ), .feedback_3_5(
        \feedback_1[7] ), .feedback_3_6(\feedback_2[8] ), 
        .feedback_3_3(\feedback_3[5] ), .feedback_3_1(\feedback_1[3] ), 
        .feedback_3_7(\feedback_2[9] ), .feedback_3_4(\feedback_0[6] ), 
        .feedback_3_0(\feedback_3[2] ), .feedback_3_2(\feedback_4[4] ), 
        .feedback_3_23(\feedback_0[25] ), .feedback_3_8(\feedback[10] )
        , .feedback_3_9(\feedback[11] ), .crc_poly_out_9(
        crc_poly_out[9]), .crc_poly_out_0(crc_poly_out[0]), 
        .crc_poly_out_4(crc_poly_out[4]), .crc_poly_out_2(
        crc_poly_out[2]), .crc_poly_out_7(crc_poly_out[7]), 
        .crc_poly_out_5(crc_poly_out[5]), .crc_poly_out_6(
        crc_poly_out[6]), .crc_poly_out_14(crc_poly_out[14]), 
        .crc_poly_out_3(crc_poly_out[3]), .crc_poly_out_11(
        crc_poly_out[11]), .feedback_5_5(\feedback_2[7] ), 
        .feedback_5_1(\feedback_3[3] ), .feedback_5_14(
        \feedback_6[16] ), .feedback_5_0(\feedback_4[2] ), 
        .feedback_5_6(\feedback[8] ), .feedback_5_2(\feedback[4] ), 
        .N_170_0(N_170_0), .N_170_0_0(N_170_0_3), .N_170_1(N_170_2), 
        .N_170_2(N_170_1), .crc_poly_size_74_0(crc_poly_size_74_0), 
        .N_170_0_1(N_170_0_6), .N_170_0_2(N_170_0_5), .N_170_0_3(
        N_170_0_4), .N_170_3(N_170), .crc_poly_size_76_0(
        crc_poly_size_76_0), .crc_poly_size_77(crc_poly_size_77), 
        .N_170_0_4(N_170_0_0), .N_170_4(N_170_4), .N_170_5(N_170_3), 
        .N_170_6(N_170_5), .N_170_0_5(N_170_0_2), .N_170_0_6(N_170_0_1)
        , .crc_poly_size_76_1(crc_poly_size_76_1), .crc_poly_size_75_0(
        crc_poly_size_75_0));
    AO1 \crc_out_1[13]  (.A(\crc_comb_out[8][13] ), .B(
        crc_poly_size_77), .C(\un65_crc_out[29]_net_1 ), .Y(
        crc_unit_out[13]));
    NOR2B \crc_out_1_RNO[15]  (.A(\crc_comb_out[8][31] ), .B(
        crc_poly_size_76_1), .Y(\un75_crc_out[31] ));
    OR3 \crc_out_1[0]  (.A(\un1_crc_out[16] ), .B(
        \crc_out_1_0[0]_net_1 ), .C(\un1_crc_out[25] ), .Y(
        crc_unit_out[0]));
    XA1 \genblk2[0].un1_crc_out[16]  (.A(\feedback[16] ), .B(
        \crc_in_masked[15] ), .C(crc_poly_size_76_0), .Y(
        \un1_crc_out[16] ));
    NOR2B \un94_poly_mux[3]  (.A(crc_poly_out[3]), .B(crc_poly_size_76)
        , .Y(\un94_poly_mux[3]_net_1 ));
    NOR2B \genblk3[31].un1_crc_init_justified[6]  (.A(crc_init_mux[6]), 
        .B(crc_poly_size_74), .Y(\un1_crc_init_justified[6] ));
    NOR2B \un105_crc_init_justified[10]  (.A(crc_init_mux[10]), .B(
        crc_poly_size_77), .Y(\un105_crc_init_justified[10]_net_1 ));
    NOR2B \un75_crc_init_justified[16]  (.A(crc_init_mux[16]), .B(
        crc_poly_size_77), .Y(\un75_crc_init_justified[16]_net_1 ));
    XA1 \un125_crc_out[25]  (.A(\feedback[25] ), .B(
        \crc_in_masked[24] ), .C(crc_poly_size_77), .Y(
        crc_unit_out[25]));
    OR2 \crc_out_1_1[1]  (.A(\un5_crc_out[25] ), .B(\crc_out_1_0[1] ), 
        .Y(\crc_out_1_1[1]_net_1 ));
    NOR2B \un35_crc_init_justified[8]  (.A(crc_init_mux[8]), .B(
        crc_poly_size_76), .Y(\un35_crc_init_justified[8]_net_1 ));
    \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_2  
        \genblk4[3].CRC_COMB  (.un100_crc_init_justified({
        \un100_crc_init_justified[11]_net_1 }), .crc_out_1_2_8(
        \crc_out_1_2[23] ), .un60_crc_init_justified_0(
        \un60_crc_init_justified[3]_net_1 ), 
        .un60_crc_init_justified_16(
        \un60_crc_init_justified[19]_net_1 ), .un15_crc_init_justified({
        \un15_crc_init_justified[28]_net_1 }), .crc_init_justified_1({
        \crc_init_justified_1[28]_net_1 }), .crc_data_in({
        crc_data_in[4]}), .crc_in_masked({\crc_in_masked_0[15] }), 
        .crc_out_1_1({\crc_out_1_1[15] }), .un104_poly_mux_16(
        \un104_poly_mux[21]_net_1 ), .un104_poly_mux_0(
        \un104_poly_mux[5]_net_1 ), .un109_poly_mux_16(
        \un109_poly_mux[22]_net_1 ), .un109_poly_mux_0(
        \un109_poly_mux[6]_net_1 ), .un79_poly_mux_16(
        \un79_poly_mux[16]_net_1 ), .un79_poly_mux_0(
        \un79_poly_mux[0]_net_1 ), .un84_poly_mux_16(
        \un84_poly_mux[17]_net_1 ), .un84_poly_mux_0(
        \un84_poly_mux[1]_net_1 ), .un89_poly_mux_16(
        \un89_poly_mux[18]_net_1 ), .un89_poly_mux_0(
        \un89_poly_mux[2]_net_1 ), .un94_poly_mux_16(
        \un94_poly_mux[19]_net_1 ), .un94_poly_mux_0(
        \un94_poly_mux[3]_net_1 ), .un99_poly_mux_16(
        \un99_poly_mux[20]_net_1 ), .un99_poly_mux_0(
        \un99_poly_mux[4]_net_1 ), .feedback_0_18(\feedback_2[31] ), 
        .feedback_0_8(\feedback_3[21] ), .feedback_0_9(
        \feedback_3[22] ), .feedback_0_7(\feedback_3[20] ), 
        .feedback_0_0(\feedback_2[13] ), .feedback_0_1(
        \feedback_2[14] ), .feedback_30(\feedback_1[31] ), 
        .feedback_12(\feedback_0[13] ), .feedback_13(\feedback_1[14] ), 
        .feedback_20(\feedback_1[21] ), .feedback_21(\feedback_2[22] ), 
        .feedback_19(\feedback_0[20] ), .feedback_14(\feedback[15] ), 
        .feedback_24(\feedback_1[25] ), .feedback_15(\feedback_3[16] ), 
        .feedback_16(\feedback_2[17] ), .feedback_17(\feedback_3[18] ), 
        .feedback_18(\feedback_2[19] ), .feedback_11(\feedback_1[12] ), 
        .feedback_5(\feedback_1[6] ), .feedback_2(\feedback_2[3] ), 
        .feedback_0_d0(\feedback[1] ), .feedback_4(\feedback_2[5] ), 
        .feedback_3(\feedback_2[4] ), .feedback_9(\feedback_2[10] ), 
        .feedback_10(\feedback_3[11] ), .feedback_7(\feedback_2[8] ), 
        .feedback_22(\feedback[23] ), .feedback_6(\feedback_2[7] ), 
        .\crc_comb_out[3] ({\crc_comb_out[3][23] }), .poly_mux_6(
        \poly_mux[12] ), .poly_mux_24(\poly_mux[30]_net_1 ), 
        .poly_mux_23(\poly_mux[29]_net_1 ), .poly_mux_9(\poly_mux[15] )
        , .poly_mux_25(\poly_mux[31]_net_1 ), .poly_mux_19(
        \poly_mux[25]_net_1 ), .poly_mux_7(\poly_mux[13] ), 
        .poly_mux_0(\poly_mux[6] ), .poly_mux_17(\poly_mux[23]_net_1 ), 
        .poly_mux_18(\poly_mux[24]_net_1 ), .\crc_comb_out[4]_15 (
        \crc_comb_out[4][15] ), .\crc_comb_out[4]_24 (
        \crc_comb_out[4][24] ), .\crc_comb_out[4]_0 (
        \crc_comb_out[4][0] ), .crc_poly_out_14(crc_poly_out[14]), 
        .crc_poly_out_3(crc_poly_out[3]), .crc_poly_out_1(
        crc_poly_out[1]), .crc_poly_out_5(crc_poly_out[5]), 
        .crc_poly_out_4(crc_poly_out[4]), .crc_poly_out_10(
        crc_poly_out[10]), .crc_poly_out_11(crc_poly_out[11]), 
        .crc_poly_out_8(crc_poly_out[8]), .crc_poly_out_7(
        crc_poly_out[7]), .crc_poly_out_0(crc_poly_out[0]), .N_170_0(
        N_170_0_3), .N_170_0_0(N_170_0_0), .N_170(N_170_1), .N_170_1(
        N_170), .N_170_2(N_170_3), .crc_poly_size_76_0(
        crc_poly_size_76_0), .crc_poly_size_77(crc_poly_size_77), 
        .crc_poly_size_75_0(crc_poly_size_75_0));
    AO1 \crc_out_1_0[2]  (.A(\crc_comb_out[8][2] ), .B(
        crc_poly_size_77), .C(\un10_crc_out[18]_net_1 ), .Y(
        \crc_out_1_0[2]_net_1 ));
    NOR2B \un25_crc_init_justified[2]  (.A(crc_init_mux[2]), .B(
        crc_poly_size_75), .Y(\un25_crc_init_justified[2]_net_1 ));
    OR2 \crc_out_1[15]  (.A(\un75_crc_out[31] ), .B(
        \un75_crc_out[15]_net_1 ), .Y(crc_unit_out[15]));
    NOR2B \un25_crc_init_justified[10]  (.A(crc_init_mux[10]), .B(
        crc_poly_size_76), .Y(\un25_crc_init_justified[10]_net_1 ));
    AO1 \crc_out_1[14]  (.A(\crc_comb_out[8][14] ), .B(
        crc_poly_size_77), .C(\un70_crc_out[30]_net_1 ), .Y(
        crc_unit_out[14]));
    NOR2B \un144_poly_mux[29]  (.A(crc_poly_out[29]), .B(
        crc_poly_size_77), .Y(\un144_poly_mux[29]_net_1 ));
    AND2 \un75_crc_out[15]  (.A(crc_poly_size_77), .B(
        \crc_comb_out[8][15] ), .Y(\un75_crc_out[15]_net_1 ));
    OR3 \crc_init_justified[24]  (.A(
        \un35_crc_init_justified[8]_net_1 ), .B(
        \un35_crc_init_justified[0]_net_1 ), .C(
        \un35_crc_init_justified[24]_net_1 ), .Y(
        \crc_init_justified[24]_net_1 ));
    NOR2B \un35_crc_out[7]  (.A(\crc_comb_out[8][7] ), .B(
        crc_poly_size_77), .Y(\un35_crc_out[7]_net_1 ));
    NOR2B \un124_poly_mux[9]  (.A(crc_poly_out[9]), .B(
        crc_poly_size_76_1), .Y(\un124_poly_mux[9]_net_1 ));
    OR3 \crc_out_1[2]  (.A(\un10_crc_out[26]_net_1 ), .B(
        \crc_out_1_0[2]_net_1 ), .C(\un10_crc_out[27]_net_1 ), .Y(
        crc_unit_out[2]));
    NOR2B \un90_crc_init_justified[13]  (.A(crc_init_mux[13]), .B(
        crc_poly_size_77), .Y(\un90_crc_init_justified[13]_net_1 ));
    NOR2B \un4_poly_mux[1]  (.A(crc_poly_out[1]), .B(crc_poly_size_77), 
        .Y(\poly_mux[1] ));
    NOR2B \un64_poly_mux[13]  (.A(crc_poly_out[13]), .B(
        crc_poly_size_77), .Y(\poly_mux[13] ));
    NOR2B \un35_crc_init_justified[24]  (.A(crc_init_mux[24]), .B(
        crc_poly_size_77), .Y(\un35_crc_init_justified[24]_net_1 ));
    AO1 \crc_out_1_1[5]  (.A(\crc_comb_out[8][29] ), .B(
        crc_poly_size_75_0), .C(\crc_out_1_0[5]_net_1 ), .Y(
        \crc_out_1_1[5]_net_1 ));
    NOR2B \un30_crc_init_justified[25]  (.A(crc_init_mux[25]), .B(
        crc_poly_size_77), .Y(\un30_crc_init_justified[25]_net_1 ));
    OR2 \poly_mux[23]  (.A(\un114_poly_mux[7]_net_1 ), .B(
        \un114_poly_mux[23]_net_1 ), .Y(\poly_mux[23]_net_1 ));
    NOR2B \un79_poly_mux[0]  (.A(crc_poly_out[0]), .B(crc_poly_size_76)
        , .Y(\un79_poly_mux[0]_net_1 ));
    NOR2B \un150_crc_out[30]  (.A(\crc_comb_out[8][30] ), .B(
        crc_poly_size_77), .Y(crc_unit_out[30]));
    NOR2B \un129_poly_mux[2]  (.A(crc_poly_out[2]), .B(
        crc_poly_size_75), .Y(\un129_poly_mux[2]_net_1 ));
    NOR2B \un70_crc_init_justified[1]  (.A(crc_init_mux[1]), .B(
        crc_poly_size_76_1), .Y(\un70_crc_init_justified[1]_net_1 ));
    NOR2B \un10_crc_init_justified[4]  (.A(crc_init_mux[4]), .B(
        crc_poly_size_74), .Y(\un10_crc_init_justified[4]_net_1 ));
    NOR2B \crc_init_justified_0_RNO[28]  (.A(crc_init_mux[4]), .B(
        crc_poly_size_75), .Y(\un15_crc_init_justified[4] ));
    NOR2B \un45_crc_init_justified[22]  (.A(crc_init_mux[22]), .B(
        crc_poly_size_77), .Y(\un45_crc_init_justified[22]_net_1 ));
    NOR2B \un134_poly_mux[27]  (.A(crc_poly_out[27]), .B(
        crc_poly_size_77), .Y(\un134_poly_mux[27]_net_1 ));
    NOR2B \un89_poly_mux[18]  (.A(crc_poly_out[18]), .B(
        crc_poly_size_77), .Y(\un89_poly_mux[18]_net_1 ));
    NOR2B \un70_crc_init_justified[17]  (.A(crc_init_mux[17]), .B(
        crc_poly_size_77), .Y(\un70_crc_init_justified[17]_net_1 ));
    NOR2B \un99_poly_mux[20]  (.A(crc_poly_out[20]), .B(
        crc_poly_size_77), .Y(\un99_poly_mux[20]_net_1 ));
    NOR2B \un30_crc_init_justified[9]  (.A(crc_init_mux[9]), .B(
        crc_poly_size_76_1), .Y(\un30_crc_init_justified[9]_net_1 ));
    NOR2B \crc_init_justified_0_RNO[27]  (.A(crc_init_mux[3]), .B(
        crc_poly_size_75_0), .Y(\un20_crc_init_justified[3] ));
    AO1 \crc_init_justified_0[29]  (.A(crc_init_mux[5]), .B(
        crc_poly_size_75_0), .C(\un10_crc_init_justified[4]_net_1 ), 
        .Y(\crc_init_justified_0[29]_net_1 ));
    NOR2B \un5_crc_init_justified[6]  (.A(crc_init_mux[6]), .B(
        crc_poly_size_75), .Y(\un5_crc_init_justified[6]_net_1 ));
    AO1 \crc_init_justified[23]  (.A(crc_init_mux[7]), .B(
        crc_poly_size_76_0), .C(\un40_crc_init_justified[23]_net_1 ), 
        .Y(\crc_init_justified[23]_net_1 ));
    \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_5  
        \genblk4[6].CRC_COMB  (.crc_out_1_5({\crc_out_1_5[15] }), 
        .un115_crc_init_justified({\un115_crc_init_justified[8]_net_1 })
        , .un75_crc_init_justified_16(
        \un75_crc_init_justified[16]_net_1 ), 
        .un75_crc_init_justified_0(\un75_crc_init_justified[0]_net_1 ), 
        .un30_crc_init_justified({\un30_crc_init_justified[25]_net_1 })
        , .crc_init_justified_1({\crc_init_justified_1[25]_net_1 }), 
        .crc_data_in({crc_data_in[1]}), .\crc_comb_out[7]_0 (
        \crc_comb_out[7][0] ), .\crc_comb_out[7]_23 (
        \crc_comb_out[7][23] ), .crc_out_1_4_0({\crc_out_1_4[23] }), 
        .un104_poly_mux_16(\un104_poly_mux[21]_net_1 ), 
        .un104_poly_mux_0(\un104_poly_mux[5]_net_1 ), 
        .un109_poly_mux_16(\un109_poly_mux[22]_net_1 ), 
        .un109_poly_mux_0(\un109_poly_mux[6]_net_1 ), 
        .un84_poly_mux_16(\un84_poly_mux[17]_net_1 ), .un84_poly_mux_0(
        \un84_poly_mux[1]_net_1 ), .un94_poly_mux_16(
        \un94_poly_mux[19]_net_1 ), .un94_poly_mux_0(
        \un94_poly_mux[3]_net_1 ), .un99_poly_mux_16(
        \un99_poly_mux[20]_net_1 ), .un99_poly_mux_0(
        \un99_poly_mux[4]_net_1 ), .un79_poly_mux_16(
        \un79_poly_mux[16]_net_1 ), .un79_poly_mux_0(
        \un79_poly_mux[0]_net_1 ), .crc_in_masked_8(
        \crc_in_masked_0[23] ), .crc_in_masked_0(\crc_in_masked_2[15] )
        , .crc_out_1_4_0_d0(\crc_out_1_4[15] ), .un89_poly_mux_16(
        \un89_poly_mux[18]_net_1 ), .un89_poly_mux_0(
        \un89_poly_mux[2]_net_1 ), .feedback_0_14(\feedback_0[23] ), 
        .feedback_0_22(\feedback_5[31] ), .feedback_0_12(
        \feedback_6[21] ), .feedback_0_13(\feedback_6[22] ), 
        .feedback_0_8(\feedback_5[17] ), .feedback_0_10(
        \feedback_5[19] ), .feedback_0_11(\feedback_6[20] ), 
        .feedback_0_5(\feedback_5[14] ), .feedback_0_0(\feedback_3[9] )
        , .feedback_0_3(\feedback_4[12] ), .feedback_0_4(
        \feedback_5[13] ), .feedback_0_6(\feedback_1[15] ), 
        .feedback_0_2(\feedback_6[11] ), .feedback_0_9(
        \feedback_6[18] ), .feedback_0_1(\feedback_4[10] ), 
        .poly_mux_29(\poly_mux[30]_net_1 ), .poly_mux_28(
        \poly_mux[29]_net_1 ), .poly_mux_27(\poly_mux[28]_net_1 ), 
        .poly_mux_26(\poly_mux[27]_net_1 ), .poly_mux_25(
        \poly_mux[26]_net_1 ), .poly_mux_30(\poly_mux[31]_net_1 ), 
        .poly_mux_23(\poly_mux[24]_net_1 ), .poly_mux_24(
        \poly_mux[25]_net_1 ), .poly_mux_14(\poly_mux[15] ), 
        .poly_mux_7(\poly_mux[8] ), .poly_mux_8(\poly_mux[9] ), 
        .poly_mux_0(\poly_mux[1] ), .poly_mux_5(\poly_mux[6] ), 
        .poly_mux_11(\poly_mux[12] ), .poly_mux_22(
        \poly_mux[23]_net_1 ), .poly_mux_12(\poly_mux[13] ), 
        .poly_mux_9(\poly_mux[10] ), .feedback_30(\feedback_4[31] ), 
        .feedback_12(\feedback_3[13] ), .feedback_13(\feedback_4[14] ), 
        .feedback_10(\feedback_2[11] ), .feedback_11(\feedback_1[12] ), 
        .feedback_8(\feedback[9] ), .feedback_9(\feedback_0[10] ), 
        .feedback_19(\feedback_3[20] ), .feedback_20(\feedback_4[21] ), 
        .feedback_17(\feedback_1[18] ), .feedback_18(\feedback_1[19] ), 
        .feedback_16(\feedback[17] ), .feedback_21(\feedback_5[22] ), 
        .feedback_25(\feedback_0[26] ), .feedback_27(\feedback_0[28] ), 
        .feedback_29(\feedback[30] ), .feedback_23(\feedback_3[24] ), 
        .feedback_24(\feedback_4[25] ), .feedback_14(\feedback_2[15] ), 
        .feedback_7(\feedback_5[8] ), .feedback_0_d0(\feedback_0[1] ), 
        .feedback_5(\feedback_4[6] ), .feedback_3(\feedback_5[4] ), 
        .feedback_4(\feedback_5[5] ), .feedback_6(\feedback_5[7] ), 
        .feedback_15(\feedback_6[16] ), .feedback_1(\feedback_4[2] ), 
        .feedback_2(\feedback_5[3] ), .crc_poly_out_0(crc_poly_out[0]), 
        .crc_poly_out_14(crc_poly_out[14]), .crc_poly_out_4(
        crc_poly_out[4]), .crc_poly_out_5(crc_poly_out[5]), 
        .crc_poly_out_7(crc_poly_out[7]), .crc_poly_out_11(
        crc_poly_out[11]), .crc_poly_out_2(crc_poly_out[2]), 
        .crc_poly_out_3(crc_poly_out[3]), .N_170_0(N_170_0_6), .N_170(
        N_170_4), .N_170_0_0(N_170_0_3), .N_170_1(N_170_2), .N_170_2(
        N_170_1), .N_170_3(N_170), .crc_poly_size_75_0(
        crc_poly_size_75_0), .crc_poly_size_77(crc_poly_size_77), 
        .crc_poly_size_76_0(crc_poly_size_76_0));
    NOR2B \un65_crc_out[29]  (.A(\crc_comb_out[8][29] ), .B(
        crc_poly_size_76_1), .Y(\un65_crc_out[29]_net_1 ));
    NOR2B \un95_crc_out[19]  (.A(\crc_comb_out[8][19] ), .B(
        crc_poly_size_77), .Y(crc_unit_out[19]));
    OR2 \crc_out_1[1]  (.A(\un5_crc_out[26]_net_1 ), .B(
        \crc_out_1_1[1]_net_1 ), .Y(crc_unit_out[1]));
    NOR2B \un55_crc_init_justified[20]  (.A(crc_init_mux[20]), .B(
        crc_poly_size_77), .Y(\un55_crc_init_justified[20]_net_1 ));
    NOR2B \un60_crc_init_justified[19]  (.A(crc_init_mux[19]), .B(
        crc_poly_size_77), .Y(\un60_crc_init_justified[19]_net_1 ));
    NOR2B \un145_crc_out[29]  (.A(\crc_comb_out[8][29] ), .B(
        crc_poly_size_77), .Y(crc_unit_out[29]));
    NOR2B \un129_poly_mux[10]  (.A(crc_poly_out[10]), .B(
        crc_poly_size_76), .Y(\un129_poly_mux[10]_net_1 ));
    NOR2B \un110_crc_init_justified[9]  (.A(crc_init_mux[9]), .B(
        crc_poly_size_77), .Y(\un110_crc_init_justified[9]_net_1 ));
    XA1 \un50_crc_out[10]  (.A(\feedback[10] ), .B(\crc_out_1_6[10] ), 
        .C(crc_poly_size_77), .Y(\un50_crc_out[10]_net_1 ));
    NOR2B \un49_poly_mux[10]  (.A(crc_poly_out[10]), .B(
        crc_poly_size_77), .Y(\poly_mux[10] ));
    OR2 \poly_mux[25]  (.A(\poly_mux_1[25]_net_1 ), .B(
        \un124_poly_mux[25]_net_1 ), .Y(\poly_mux[25]_net_1 ));
    XA1 \un80_crc_out[16]  (.A(\feedback[16] ), .B(\crc_in_masked[15] )
        , .C(crc_poly_size_77), .Y(crc_unit_out[16]));
    NOR2B \un124_poly_mux[0]  (.A(crc_poly_out[0]), .B(
        crc_poly_size_74), .Y(\un124_poly_mux[0]_net_1 ));
    AND2 \un20_crc_init_justified[11]  (.A(crc_poly_size_76), .B(
        crc_init_mux[11]), .Y(\un20_crc_init_justified[11]_net_1 ));
    AO1 \crc_out_1_0[6]  (.A(\crc_comb_out[8][6] ), .B(
        crc_poly_size_77), .C(\un30_crc_out[22]_net_1 ), .Y(
        \crc_out_1_0[6]_net_1 ));
    AO1 \crc_init_justified_1[29]  (.A(crc_init_mux[13]), .B(
        crc_poly_size_76_0), .C(\crc_init_justified_0[29]_net_1 ), .Y(
        \crc_init_justified_1[29]_net_1 ));
    NOR2B \un60_crc_init_justified[3]  (.A(crc_init_mux[3]), .B(
        crc_poly_size_76), .Y(\un60_crc_init_justified[3]_net_1 ));
    AND2 \un5_crc_out[1]  (.A(crc_poly_size_77), .B(
        \crc_comb_out[8][1] ), .Y(\un5_crc_out[1]_net_1 ));
    NOR2B \un134_poly_mux[11]  (.A(crc_poly_out[11]), .B(
        crc_poly_size_76), .Y(\un134_poly_mux[11]_net_1 ));
    NOR2B \un109_poly_mux[22]  (.A(crc_poly_out[22]), .B(
        crc_poly_size_77), .Y(\un109_poly_mux[22]_net_1 ));
    AO1 \crc_init_justified[21]  (.A(crc_init_mux[5]), .B(
        crc_poly_size_76_0), .C(\un50_crc_init_justified[21]_net_1 ), 
        .Y(\crc_init_justified[21]_net_1 ));
    NOR2B \un124_poly_mux[1]  (.A(crc_poly_out[1]), .B(
        crc_poly_size_75), .Y(\un124_poly_mux[1]_net_1 ));
    NOR2B \un65_crc_init_justified[2]  (.A(crc_init_mux[2]), .B(
        crc_poly_size_76_1), .Y(\un65_crc_init_justified[2]_net_1 ));
    OR3 \crc_out_1[6]  (.A(\un30_crc_out[31]_net_1 ), .B(
        \crc_out_1_0[6]_net_1 ), .C(\un30_crc_out[30]_net_1 ), .Y(
        crc_unit_out[6]));
    OR3 \poly_mux_1[30]  (.A(\un149_poly_mux[6]_net_1 ), .B(
        \un149_poly_mux[5]_net_1 ), .C(\un149_poly_mux[14]_net_1 ), .Y(
        \poly_mux_1[30]_net_1 ));
    NOR2B \un5_crc_init_justified[5]  (.A(crc_init_mux[5]), .B(
        crc_poly_size_74), .Y(\un5_crc_init_justified[5]_net_1 ));
    AO1 \crc_out_1[8]  (.A(\crc_comb_out[8][24] ), .B(
        crc_poly_size_76_0), .C(\un40_crc_out[8]_net_1 ), .Y(
        crc_unit_out[8]));
    NOR2B \un29_poly_mux[6]  (.A(crc_poly_out[6]), .B(crc_poly_size_77)
        , .Y(\poly_mux[6] ));
    NOR2B \un15_crc_out[19]  (.A(\crc_comb_out[8][19] ), .B(
        crc_poly_size_76), .Y(\un15_crc_out[19]_net_1 ));
    NOR2B \un149_poly_mux[5]  (.A(crc_poly_out[5]), .B(
        crc_poly_size_74), .Y(\un149_poly_mux[5]_net_1 ));
    NOR2B \un85_crc_init_justified[14]  (.A(crc_init_mux[14]), .B(
        crc_poly_size_77), .Y(\un85_crc_init_justified[14]_net_1 ));
    NOR2B \un109_poly_mux[6]  (.A(crc_poly_out[6]), .B(
        crc_poly_size_76), .Y(\un109_poly_mux[6]_net_1 ));
    \crc_comb_32s_4294967295_genblk4[0].CRC_COMB_1  
        \genblk4[2].CRC_COMB  (.\crc_comb_out[2] ({
        \crc_comb_out[2][23] }), .crc_out_1_1({\crc_out_1_1[15] }), 
        .un95_crc_init_justified({\un95_crc_init_justified[12]_net_1 })
        , .un55_crc_init_justified_16(
        \un55_crc_init_justified[20]_net_1 ), 
        .un55_crc_init_justified_0(\un55_crc_init_justified[4]_net_1 ), 
        .un10_crc_init_justified({\un10_crc_init_justified[29]_net_1 })
        , .crc_init_justified_1({\crc_init_justified_1[29]_net_1 }), 
        .crc_data_in({crc_data_in[5]}), .\crc_comb_out[3] ({
        \crc_comb_out[3][24] , \crc_comb_out[3][23] }), 
        .crc_in_masked_1(\crc_in_masked_1[24] ), .crc_out_1_0_1(
        \crc_out_1_0[24] ), .un104_poly_mux_16(
        \un104_poly_mux[21]_net_1 ), .un104_poly_mux_0(
        \un104_poly_mux[5]_net_1 ), .un79_poly_mux_16(
        \un79_poly_mux[16]_net_1 ), .un79_poly_mux_0(
        \un79_poly_mux[0]_net_1 ), .un84_poly_mux_16(
        \un84_poly_mux[17]_net_1 ), .un84_poly_mux_0(
        \un84_poly_mux[1]_net_1 ), .un89_poly_mux_16(
        \un89_poly_mux[18]_net_1 ), .un89_poly_mux_0(
        \un89_poly_mux[2]_net_1 ), .un94_poly_mux_16(
        \un94_poly_mux[19]_net_1 ), .un94_poly_mux_0(
        \un94_poly_mux[3]_net_1 ), .un99_poly_mux_16(
        \un99_poly_mux[20]_net_1 ), .un99_poly_mux_0(
        \un99_poly_mux[4]_net_1 ), .crc_poly_out_9(crc_poly_out[11]), 
        .crc_poly_out_3(crc_poly_out[5]), .crc_poly_out_0(
        crc_poly_out[2]), .crc_poly_out_2(crc_poly_out[4]), 
        .crc_poly_out_1(crc_poly_out[3]), .crc_poly_out_5(
        crc_poly_out[7]), .crc_poly_out_12(crc_poly_out[14]), 
        .feedback_0_11(\feedback_1[24] ), .feedback_0_18(
        \feedback_1[31] ), .feedback_0_8(\feedback_2[21] ), 
        .feedback_0_0(\feedback_1[13] ), .feedback_0_1(
        \feedback_1[14] ), .feedback_0_9(\feedback_2[22] ), 
        .un109_poly_mux_16(\un109_poly_mux[22]_net_1 ), 
        .un109_poly_mux_0(\un109_poly_mux[6]_net_1 ), .feedback_29(
        \feedback_0[31] ), .feedback_11(\feedback[13] ), .feedback_12(
        \feedback_0[14] ), .feedback_19(\feedback_0[21] ), 
        .feedback_20(\feedback_1[22] ), .feedback_14(\feedback_2[16] ), 
        .feedback_15(\feedback_1[17] ), .feedback_16(\feedback_2[18] ), 
        .feedback_17(\feedback_1[19] ), .feedback_18(\feedback_2[20] ), 
        .feedback_9(\feedback_2[11] ), .feedback_10(\feedback_0[12] ), 
        .feedback_13(\feedback[15] ), .feedback_6(\feedback_1[8] ), 
        .feedback_3(\feedback_1[5] ), .feedback_0_d0(\feedback_1[2] ), 
        .feedback_2(\feedback_1[4] ), .feedback_1(\feedback_1[3] ), 
        .feedback_7(\feedback_0[9] ), .feedback_8(\feedback_1[10] ), 
        .feedback_5(\feedback_1[7] ), .feedback_4(\feedback_0[6] ), 
        .poly_mux_18(\poly_mux[24]_net_1 ), .poly_mux_24(
        \poly_mux[30]_net_1 ), .poly_mux_25(\poly_mux[31]_net_1 ), 
        .poly_mux_6(\poly_mux[12] ), .poly_mux_7(\poly_mux[13] ), 
        .poly_mux_9(\poly_mux[15] ), .poly_mux_2(\poly_mux[8] ), 
        .poly_mux_3(\poly_mux[9] ), .poly_mux_4(\poly_mux[10] ), 
        .poly_mux_0(\poly_mux[6] ), .poly_mux_17(\poly_mux[23]_net_1 ), 
        .N_170_0(N_170_0_2), .crc_poly_size_75(crc_poly_size_75), 
        .N_170(N_170_2), .N_170_0_0(N_170_0_0), .crc_poly_size_74_0(
        crc_poly_size_74_0), .crc_poly_size_77(crc_poly_size_77));
    NOR2B \un15_crc_init_justified[28]  (.A(crc_init_mux[28]), .B(
        crc_poly_size_77), .Y(\un15_crc_init_justified[28]_net_1 ));
    NOR2B \un55_crc_init_justified[4]  (.A(crc_init_mux[4]), .B(
        crc_poly_size_76_1), .Y(\un55_crc_init_justified[4]_net_1 ));
    NOR2B \un80_crc_init_justified[15]  (.A(crc_init_mux[15]), .B(
        crc_poly_size_77), .Y(\un80_crc_init_justified[15]_net_1 ));
    AND2 \un15_crc_init_justified[12]  (.A(crc_poly_size_76), .B(
        crc_init_mux[12]), .Y(\un15_crc_init_justified[12]_net_1 ));
    NOR2B \un149_poly_mux[14]  (.A(crc_poly_out[14]), .B(
        crc_poly_size_76), .Y(\un149_poly_mux[14]_net_1 ));
    NOR2B \un50_crc_init_justified[21]  (.A(crc_init_mux[21]), .B(
        crc_poly_size_77), .Y(\un50_crc_init_justified[21]_net_1 ));
    NOR2B \un124_poly_mux[25]  (.A(crc_poly_out[25]), .B(
        crc_poly_size_77), .Y(\un124_poly_mux[25]_net_1 ));
    NOR2B \un35_crc_init_justified[0]  (.A(crc_init_mux[0]), .B(
        crc_poly_size_75), .Y(\un35_crc_init_justified[0]_net_1 ));
    OR3 \crc_init_justified_1[25]  (.A(
        \un30_crc_init_justified[1]_net_1 ), .B(
        \un30_crc_init_justified[0]_net_1 ), .C(
        \un30_crc_init_justified[9]_net_1 ), .Y(
        \crc_init_justified_1[25]_net_1 ));
    NOR2B \un119_poly_mux[24]  (.A(crc_poly_out[24]), .B(
        crc_poly_size_77), .Y(\un119_poly_mux[24]_net_1 ));
    AO1 \crc_init_justified[31]  (.A(crc_init_mux[31]), .B(
        crc_poly_size_77), .C(\crc_init_justified_1[31]_net_1 ), .Y(
        \crc_init_justified[31]_net_1 ));
    OR3 \poly_mux[29]  (.A(\poly_mux_0[29]_net_1 ), .B(
        \un144_poly_mux[13]_net_1 ), .C(\un144_poly_mux[29]_net_1 ), 
        .Y(\poly_mux[29]_net_1 ));
    NOR2B \un74_poly_mux[15]  (.A(crc_poly_out[15]), .B(
        crc_poly_size_77), .Y(\poly_mux[15] ));
    XA1 \un55_crc_out[11]  (.A(\feedback[11] ), .B(\crc_out_1_6[11] ), 
        .C(crc_poly_size_77), .Y(\un55_crc_out[11]_net_1 ));
    NOR2B \un25_crc_init_justified[26]  (.A(crc_init_mux[26]), .B(
        crc_poly_size_77), .Y(\un25_crc_init_justified[26]_net_1 ));
    NOR2B \un130_crc_out[26]  (.A(\crc_comb_out[8][26] ), .B(
        crc_poly_size_77), .Y(crc_unit_out[26]));
    AO1 \crc_out_1[7]  (.A(\crc_comb_out[8][31] ), .B(
        crc_poly_size_75_0), .C(\crc_out_1_0[7]_net_1 ), .Y(
        crc_unit_out[7]));
    NOR2B \un89_poly_mux[2]  (.A(crc_poly_out[2]), .B(crc_poly_size_76)
        , .Y(\un89_poly_mux[2]_net_1 ));
    NOR2B \un70_crc_out[30]  (.A(\crc_comb_out[8][30] ), .B(
        crc_poly_size_76), .Y(\un70_crc_out[30]_net_1 ));
    NOR2B \un95_crc_init_justified[12]  (.A(crc_init_mux[12]), .B(
        crc_poly_size_77), .Y(\un95_crc_init_justified[12]_net_1 ));
    NOR2B \un44_poly_mux[9]  (.A(crc_poly_out[9]), .B(crc_poly_size_77)
        , .Y(\poly_mux[9] ));
    \crc_comb_32s_4294967295_genblk4[0].CRC_COMB  
        \genblk4[0].CRC_COMB  (.crc_data_in({crc_data_in[7]}), 
        .crc_init_justified({\crc_init_justified[31]_net_1 }), 
        .un79_poly_mux_16(\un79_poly_mux[16]_net_1 ), .un79_poly_mux_0(
        \un79_poly_mux[0]_net_1 ), .un84_poly_mux_16(
        \un84_poly_mux[17]_net_1 ), .un84_poly_mux_0(
        \un84_poly_mux[1]_net_1 ), .un89_poly_mux_16(
        \un89_poly_mux[18]_net_1 ), .un89_poly_mux_0(
        \un89_poly_mux[2]_net_1 ), .un94_poly_mux_16(
        \un94_poly_mux[19]_net_1 ), .un94_poly_mux_0(
        \un94_poly_mux[3]_net_1 ), .un109_poly_mux_16(
        \un109_poly_mux[22]_net_1 ), .un109_poly_mux_0(
        \un109_poly_mux[6]_net_1 ), .un99_poly_mux_16(
        \un99_poly_mux[20]_net_1 ), .un99_poly_mux_0(
        \un99_poly_mux[4]_net_1 ), .\crc_comb_out[1] ({
        \crc_comb_out[1][0] }), .crc_poly_out_14(crc_poly_out[14]), 
        .crc_poly_out_3(crc_poly_out[3]), .crc_poly_out_11(
        crc_poly_out[11]), .crc_poly_out_0(crc_poly_out[0]), 
        .crc_poly_out_2(crc_poly_out[2]), .crc_poly_out_7(
        crc_poly_out[7]), .crc_poly_out_5(crc_poly_out[5]), 
        .poly_mux_4(\poly_mux[13] ), .poly_mux_16(\poly_mux[25]_net_1 )
        , .poly_mux_15(\poly_mux[24]_net_1 ), .poly_mux_22(
        \poly_mux[31]_net_1 ), .poly_mux_0(\poly_mux[9] ), 
        .feedback_11(\feedback[13] ), .feedback_12(\feedback[14] ), 
        .feedback_23(\feedback_0[25] ), .feedback_14(\feedback_0[16] ), 
        .feedback_15(\feedback[17] ), .feedback_22(\feedback_0[24] ), 
        .feedback_1(\feedback[3] ), .feedback_16(\feedback_0[18] ), 
        .feedback_17(\feedback[19] ), .feedback_20(\feedback_0[22] ), 
        .feedback_9(\feedback_0[11] ), .feedback_18(\feedback_0[20] ), 
        .feedback_0(\feedback[2] ), .feedback_5(\feedback[7] ), 
        .feedback_29(\feedback[31] ), .feedback_3(\feedback[5] ), 
        .feedback_7(\feedback[9] ), .feedback_19(\feedback_0[21] ), 
        .un104_poly_mux_16(\un104_poly_mux[21]_net_1 ), 
        .un104_poly_mux_0(\un104_poly_mux[5]_net_1 ), .N_170_0(
        N_170_0_0), .N_170(N_170), .crc_poly_size_77(crc_poly_size_77));
    NOR2B \un59_poly_mux[12]  (.A(crc_poly_out[12]), .B(
        crc_poly_size_77), .Y(\poly_mux[12] ));
    AO1 \crc_out_1_0[3]  (.A(\crc_comb_out[8][3] ), .B(
        crc_poly_size_77), .C(\un15_crc_out[19]_net_1 ), .Y(
        \crc_out_1_0[3]_net_1 ));
    AO1 \poly_mux_0[31]  (.A(crc_poly_out[7]), .B(crc_poly_size_75_0), 
        .C(\un154_poly_mux[6] ), .Y(\poly_mux_0[31]_net_1 ));
    AO1 \crc_out_1_0[7]  (.A(\crc_comb_out[8][23] ), .B(
        crc_poly_size_76_0), .C(\un35_crc_out[7]_net_1 ), .Y(
        \crc_out_1_0[7]_net_1 ));
    OR3 \crc_init_justified_1[26]  (.A(
        \un25_crc_init_justified[2]_net_1 ), .B(
        \un25_crc_init_justified[1]_net_1 ), .C(
        \un25_crc_init_justified[10]_net_1 ), .Y(
        \crc_init_justified_1[26]_net_1 ));
    XA1 \un105_crc_out[21]  (.A(\feedback[21] ), .B(\crc_out_1_4[21] ), 
        .C(crc_poly_size_77), .Y(crc_unit_out[21]));
    OR3 \poly_mux[31]  (.A(\poly_mux_0[31]_net_1 ), .B(
        \un154_poly_mux[15] ), .C(\un154_poly_mux[31] ), .Y(
        \poly_mux[31]_net_1 ));
    NOR2B \un30_crc_init_justified[1]  (.A(crc_init_mux[1]), .B(
        crc_poly_size_75_0), .Y(\un30_crc_init_justified[1]_net_1 ));
    XA1 \un45_crc_out[25]  (.A(\feedback[25] ), .B(\crc_in_masked[24] )
        , .C(crc_poly_size_76_1), .Y(\un45_crc_out[25]_net_1 ));
    
endmodule


module crc_datapath(
       crc_poly_size,
       state_byte_i,
       state_byte,
       state_byte_0,
       size_in,
       bus_size,
       bus_wr_0,
       bus_wr_1,
       bus_wr_16,
       bus_wr_25,
       bus_wr_2,
       bus_wr_3,
       crc_idr_out,
       crc_out,
       crc_init_out,
       crc_poly_out,
       rev_in_type_0,
       rev_in_type,
       FAB_CLK,
       N_56,
       crc_init_en,
       byte_en_0,
       byte_en,
       crc_poly_en,
       N_348,
       N_350,
       N_352,
       N_353,
       crc_poly_en_0,
       N_358,
       N_360,
       N_361,
       N_364,
       N_365,
       N_366,
       N_332,
       N_333,
       N_334,
       N_335,
       N_336,
       N_337,
       crc_idr_en,
       N_347,
       buffer_en_0,
       buffer_en,
       rev_out_type_0,
       rev_out_type,
       N_118_1,
       crc_ahb_ip_MSS_0_M2F_RESET_N,
       N_128,
       N_294_0,
       bypass_byte0,
       crc_init_en_0,
       N_367,
       crc_poly_size_77,
       N_349,
       N_357,
       N_356,
       N_354,
       N_351,
       N_362,
       N_355,
       N_363,
       crc_poly_size_77_0
    );
input  [1:0] crc_poly_size;
input  [0:0] state_byte_i;
input  [4:4] state_byte;
input  [4:4] state_byte_0;
output [1:0] size_in;
input  [1:0] bus_size;
input  bus_wr_0;
input  bus_wr_1;
input  bus_wr_16;
input  bus_wr_25;
input  bus_wr_2;
input  bus_wr_3;
output [7:0] crc_idr_out;
output [31:0] crc_out;
output [31:0] crc_init_out;
output [31:0] crc_poly_out;
input  [0:0] rev_in_type_0;
input  [1:0] rev_in_type;
input  FAB_CLK;
input  N_56;
input  crc_init_en;
input  byte_en_0;
input  byte_en;
input  crc_poly_en;
input  N_348;
input  N_350;
input  N_352;
input  N_353;
input  crc_poly_en_0;
input  N_358;
input  N_360;
input  N_361;
input  N_364;
input  N_365;
input  N_366;
input  N_332;
input  N_333;
input  N_334;
input  N_335;
input  N_336;
input  N_337;
input  crc_idr_en;
input  N_347;
input  buffer_en_0;
input  buffer_en;
input  rev_out_type_0;
input  rev_out_type;
input  N_118_1;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;
input  N_128;
input  N_294_0;
input  bypass_byte0;
input  crc_init_en_0;
input  N_367;
output crc_poly_size_77;
input  N_349;
input  N_357;
input  N_356;
input  N_354;
input  N_351;
input  N_362;
input  N_355;
input  N_363;
input  crc_poly_size_77_0;

    wire crc_init_sel_ff_0, crc_init_sel_ff_RNI2BI2B_net_1, 
        crc_poly_size_75_0_net_1, crc_poly_size_76_1_net_1, 
        crc_poly_size_76_0_net_1, crc_poly_size_74_0_net_1, 
        un1_crc_init_en_1_0_net_1, N_165, crc_init_sel_ff_net_1, N_166, 
        \byte_ff[0]_net_1 , \buffer_ff[0]_net_1 , N_167, 
        \byte_ff[1]_net_1 , \buffer_ff[1]_net_1 , N_168, 
        \byte_ff[2]_net_1 , \buffer_ff[2]_net_1 , N_169, 
        \byte_ff[3]_net_1 , \buffer_ff[3]_net_1 , N_170, 
        \byte_ff[4]_net_1 , \buffer_ff[4]_net_1 , N_171, 
        \byte_ff[5]_net_1 , \buffer_ff[5]_net_1 , N_172, 
        \byte_ff[6]_net_1 , \buffer_ff[6]_net_1 , N_173, 
        \byte_ff[7]_net_1 , \buffer_ff[7]_net_1 , N_175, 
        \byte_ff[9]_net_1 , \buffer_ff[9]_net_1 , N_176, 
        \byte_ff[10]_net_1 , \buffer_ff[10]_net_1 , N_178, 
        \byte_ff[12]_net_1 , \buffer_ff[12]_net_1 , N_179, 
        \byte_ff[13]_net_1 , \buffer_ff[13]_net_1 , N_181, 
        \byte_ff[15]_net_1 , \buffer_ff[15]_net_1 , N_182, 
        \byte_ff[16]_net_1 , \buffer_ff[16]_net_1 , N_183, 
        \byte_ff[17]_net_1 , \buffer_ff[17]_net_1 , N_184, 
        \byte_ff[18]_net_1 , \buffer_ff[18]_net_1 , N_185, 
        \byte_ff[19]_net_1 , \buffer_ff[19]_net_1 , N_187, 
        \byte_ff[21]_net_1 , \buffer_ff[21]_net_1 , N_189, 
        \byte_ff[23]_net_1 , \buffer_ff[23]_net_1 , N_190, 
        \byte_ff[24]_net_1 , \buffer_ff[24]_net_1 , N_191, 
        \byte_ff[25]_net_1 , \buffer_ff[25]_net_1 , N_192, 
        \byte_ff[26]_net_1 , \buffer_ff[26]_net_1 , N_193, 
        \byte_ff[27]_net_1 , \buffer_ff[27]_net_1 , N_194, 
        \byte_ff[28]_net_1 , \buffer_ff[28]_net_1 , N_195, 
        \byte_ff[29]_net_1 , \buffer_ff[29]_net_1 , N_197, 
        \byte_ff[31]_net_1 , \buffer_ff[31]_net_1 , N_198, N_199, 
        N_203, N_205, N_207, N_208, N_213, N_214, N_215, N_216, N_219, 
        N_220, N_221, N_223, N_224, N_225, N_226, N_227, N_228, N_229, 
        N_230, N_231, N_234, N_235, N_237, N_239, \crc_unit_out[1] , 
        \crc_out_ff[1]_net_1 , N_240, \crc_unit_out[2] , 
        \crc_out_ff[2]_net_1 , N_241, \crc_unit_out[3] , 
        \crc_out_ff[3]_net_1 , N_247, \crc_unit_out[9] , 
        \crc_out_ff[9]_net_1 , N_248, \crc_unit_out[10] , 
        \crc_out_ff[10]_net_1 , N_253, \crc_unit_out[15] , 
        \crc_out_ff[15]_net_1 , N_254, \crc_unit_out[16] , 
        \crc_out_ff[16]_net_1 , N_259, \crc_unit_out[21] , 
        \crc_out_ff[21]_net_1 , N_260, \crc_unit_out[22] , 
        \crc_out_ff[22]_net_1 , N_263, \crc_unit_out[25] , 
        \crc_out_ff[25]_net_1 , N_265, \crc_unit_out[27] , 
        \crc_out_ff[27]_net_1 , N_266, \crc_unit_out[28] , 
        \crc_out_ff[28]_net_1 , N_267, \crc_unit_out[29] , 
        \crc_out_ff[29]_net_1 , N_269, \crc_unit_out[31] , 
        \crc_out_ff[31]_net_1 , N_270, \bus_reversed[0] , N_271, 
        \bus_reversed[1] , N_272, \bus_reversed[2] , N_273, 
        \bus_reversed[3] , N_275, \bus_reversed[5] , N_276, 
        \bus_reversed[6] , N_277, \bus_reversed[7] , N_279, 
        \bus_reversed[9] , N_280, \bus_reversed[10] , N_283, 
        \bus_reversed[13] , N_285, \bus_reversed[15] , N_286, 
        \bus_reversed[16] , N_287, \bus_reversed[17] , N_288, 
        \bus_reversed[18] , N_289, \bus_reversed[19] , N_291, 
        \bus_reversed[21] , N_293, \bus_reversed[23] , N_294, 
        \bus_reversed[24] , N_295, \bus_reversed[25] , N_296, 
        \bus_reversed[26] , N_297, \bus_reversed[27] , N_298, 
        \bus_reversed[28] , N_299, \bus_reversed[29] , N_301, 
        \bus_reversed[31] , N_129, \size_ff[0]_net_1 , 
        \bf_size_ff[0]_net_1 , N_130, \size_ff[1]_net_1 , 
        \bf_size_ff[1]_net_1 , N_132, \crc_init_ff_3[1] , N_133, 
        \crc_init_ff_3[2] , N_134, \crc_init_ff_3[3] , N_135, 
        \crc_init_ff_3[4] , N_136, \crc_init_ff_3[5] , N_140, 
        \crc_init_ff_3[9] , N_141, \crc_init_ff_3[10] , N_146, 
        \crc_init_ff_3[15] , N_147, \crc_init_ff_3[16] , 
        un1_crc_init_en_1_net_1, N_148, \crc_init_ff_3[17] , N_152, 
        \crc_init_ff_3[21] , N_153, \crc_init_ff_3[22] , N_154, 
        \crc_init_ff_3[23] , N_155, \crc_init_ff_3[24] , N_156, 
        \crc_init_ff_3[25] , N_158, \crc_init_ff_3[27] , N_159, 
        \crc_init_ff_3[28] , N_160, \crc_init_ff_3[29] , N_162, 
        \crc_init_ff_3[31] , N_163, \bf_size_ff_4[0] , 
        un1_buffer_en_net_1, N_164, \bf_size_ff_4[1] , 
        \crc_init_mux[0] , \crc_out_ff[0]_net_1 , \crc_init_mux[31] , 
        \crc_out_ff[30]_net_1 , \crc_init_mux[2] , \crc_init_mux[3] , 
        \crc_init_mux[28] , \crc_init_mux[29] , \crc_init_mux[4] , 
        \crc_out_ff[4]_net_1 , \crc_init_mux[5] , 
        \crc_out_ff[5]_net_1 , \crc_init_mux[26] , 
        \crc_out_ff[26]_net_1 , \crc_init_mux[27] , \crc_init_mux[24] , 
        \crc_out_ff[24]_net_1 , \crc_init_mux[25] , 
        \crc_out_ff[7]_net_1 , \crc_out_ff[6]_net_1 , 
        \crc_init_mux[8] , \crc_out_ff[8]_net_1 , \crc_init_mux[9] , 
        \crc_init_mux[22] , \crc_out_ff[23]_net_1 , \crc_init_mux[10] , 
        \crc_init_mux[11] , \crc_out_ff[11]_net_1 , \crc_init_mux[21] , 
        \crc_init_mux[12] , \crc_out_ff[12]_net_1 , \crc_init_mux[13] , 
        \crc_out_ff[13]_net_1 , \crc_init_mux[18] , 
        \crc_out_ff[18]_net_1 , \crc_init_mux[19] , 
        \crc_out_ff[19]_net_1 , \crc_init_mux[15] , \crc_init_mux[16] , 
        \crc_init_mux[17] , \crc_out_ff[17]_net_1 , 
        \crc_out_ff[14]_net_1 , \crc_out_ff_RNO[1]_net_1 , 
        \crc_out_ff_RNO[2]_net_1 , \crc_poly_ff_RNO[5]_net_1 , 
        \crc_poly_ff_RNO[7]_net_1 , \crc_poly_ff_RNO[10]_net_1 , 
        \crc_poly_ff_RNO[16]_net_1 , \crc_poly_ff_RNO[22]_net_1 , 
        \crc_poly_ff_RNO[23]_net_1 , \crc_poly_ff_RNO[26]_net_1 , 
        \bf_size_ff_RNO[1]_net_1 , \size_ff_RNO[1]_net_1 , 
        \crc_init_ff_RNO[22]_net_1 , \crc_init_ff_RNO[23]_net_1 , 
        \crc_init_ff_RNO[24]_net_1 , \crc_init_ff_RNO[25]_net_1 , 
        \crc_init_ff_RNO[27]_net_1 , \crc_init_ff_RNO[28]_net_1 , 
        \crc_init_ff_RNO[29]_net_1 , \crc_init_ff_RNO[31]_net_1 , 
        \crc_poly_ff_RNO[0]_net_1 , \crc_poly_ff_RNO[1]_net_1 , 
        \crc_init_ff_RNO[9]_net_1 , \crc_init_ff_RNO[10]_net_1 , 
        \crc_init_ff_RNO[15]_net_1 , \crc_init_ff_RNO[16]_net_1 , 
        \crc_init_ff_RNO[17]_net_1 , \crc_init_ff_RNO[21]_net_1 , 
        \byte_ff_RNO[28]_net_1 , \byte_ff_RNO[29]_net_1 , 
        \byte_ff_RNO[31]_net_1 , \crc_init_ff_RNO[1]_net_1 , 
        \crc_init_ff_RNO[2]_net_1 , \crc_init_ff_RNO[3]_net_1 , 
        \crc_init_ff_RNO[4]_net_1 , \crc_init_ff_RNO[5]_net_1 , 
        \byte_ff_RNO[15]_net_1 , \byte_ff_RNO[16]_net_1 , 
        \byte_ff_RNO[17]_net_1 , \byte_ff_RNO[18]_net_1 , 
        \byte_ff_RNO[19]_net_1 , \byte_ff_RNO[21]_net_1 , 
        \byte_ff_RNO[23]_net_1 , \byte_ff_RNO[24]_net_1 , 
        \byte_ff_RNO[25]_net_1 , \byte_ff_RNO[26]_net_1 , 
        \byte_ff_RNO[27]_net_1 , \byte_ff_RNO[2]_net_1 , 
        \byte_ff_RNO[3]_net_1 , \byte_ff_RNO[4]_net_1 , 
        \byte_ff_RNO[5]_net_1 , \byte_ff_RNO[6]_net_1 , 
        \byte_ff_RNO[7]_net_1 , \byte_ff_RNO[9]_net_1 , 
        \byte_ff_RNO[10]_net_1 , \byte_ff_RNO[12]_net_1 , 
        \byte_ff_RNO[13]_net_1 , \buffer_ff_RNO[21]_net_1 , 
        \buffer_ff_RNO[23]_net_1 , \buffer_ff_RNO[24]_net_1 , 
        \buffer_ff_RNO[25]_net_1 , \buffer_ff_RNO[26]_net_1 , 
        \buffer_ff_RNO[27]_net_1 , \buffer_ff_RNO[28]_net_1 , 
        \buffer_ff_RNO[29]_net_1 , \buffer_ff_RNO[31]_net_1 , 
        \byte_ff_RNO[0]_net_1 , \byte_ff_RNO[1]_net_1 , 
        \buffer_ff_RNO[9]_net_1 , \buffer_ff_RNO[10]_net_1 , 
        \buffer_ff_RNO[13]_net_1 , \buffer_ff_RNO[15]_net_1 , 
        \buffer_ff_RNO[16]_net_1 , \buffer_ff_RNO[17]_net_1 , 
        \buffer_ff_RNO[18]_net_1 , \buffer_ff_RNO[19]_net_1 , 
        \crc_poly_ff_RNO[29]_net_1 , \crc_poly_ff_RNO[30]_net_1 , 
        \crc_poly_ff_RNO[31]_net_1 , \bf_size_ff_RNO[0]_net_1 , 
        \size_ff_RNO[0]_net_1 , \buffer_ff_RNO[0]_net_1 , 
        \buffer_ff_RNO[1]_net_1 , \buffer_ff_RNO[2]_net_1 , 
        \buffer_ff_RNO[3]_net_1 , \buffer_ff_RNO[5]_net_1 , 
        \buffer_ff_RNO[6]_net_1 , \buffer_ff_RNO[7]_net_1 , 
        \crc_poly_ff_RNO[9]_net_1 , \crc_poly_ff_RNO[15]_net_1 , 
        \crc_poly_ff_RNO[17]_net_1 , \crc_poly_ff_RNO[18]_net_1 , 
        \crc_poly_ff_RNO[21]_net_1 , \crc_poly_ff_RNO[25]_net_1 , 
        \crc_poly_ff_RNO[27]_net_1 , \crc_poly_ff_RNO[28]_net_1 , 
        \crc_out_ff_RNO[29]_net_1 , \crc_out_ff_RNO[31]_net_1 , 
        \crc_idr_ff_RNO[0]_net_1 , \crc_idr_ff_RNO[1]_net_1 , 
        \crc_idr_ff_RNO[4]_net_1 , \crc_idr_ff_RNO[5]_net_1 , 
        \crc_idr_ff_RNO[7]_net_1 , \crc_out_ff_RNO[16]_net_1 , 
        \crc_out_ff_RNO[21]_net_1 , \crc_out_ff_RNO[22]_net_1 , 
        \crc_out_ff_RNO[25]_net_1 , \crc_out_ff_RNO[27]_net_1 , 
        \crc_out_ff_RNO[28]_net_1 , \crc_out_ff_RNO[3]_net_1 , 
        \crc_out_ff_RNO[9]_net_1 , \crc_out_ff_RNO[10]_net_1 , 
        \crc_out_ff_RNO[15]_net_1 , N_96, \crc_data_in0[0] , N_97, 
        \crc_data_in0[1] , N_98, \crc_data_in0[2] , N_99, 
        \crc_data_in0[3] , N_100, \byte_ff[20]_net_1 , 
        \crc_data_in0[4] , N_101, \crc_data_in0[5] , N_103, 
        \crc_data_in0[7] , N_104, \byte_ff[8]_net_1 , N_105, N_106, 
        N_107, \byte_ff[11]_net_1 , N_108, N_109, N_111, 
        \crc_data_in[0] , \crc_data_in[1] , \crc_data_in[2] , 
        \crc_data_in[3] , \crc_data_in[4] , \crc_data_in[5] , 
        \crc_data_in[7] , crc_poly_size_74_net_1, 
        crc_poly_size_76_net_1, \crc_out_ff_RNO[7]_net_1 , N_245, 
        \crc_out_ff_RNO[23]_net_1 , N_261, \buffer_ff_RNO[8]_net_1 , 
        N_278, \byte_ff_RNO[8]_net_1 , N_174, \buffer_ff[8]_net_1 , 
        \bus_reversed[8] , \crc_unit_out[23] , \crc_unit_out[7] , 
        \crc_init_ff_3[6] , \crc_poly_ff_RNO[14]_net_1 , N_212, 
        \buffer_ff_RNO[14]_net_1 , N_284, \crc_init_ff_RNO[6]_net_1 , 
        N_137, \buffer_ff[14]_net_1 , \bus_reversed[14] , 
        \crc_init_ff_3[18] , \crc_init_ff_3[13] , 
        \crc_out_ff_RNO[13]_net_1 , N_251, \crc_out_ff_RNO[18]_net_1 , 
        N_256, \crc_poly_ff_RNO[13]_net_1 , N_211, 
        \crc_init_ff_RNO[18]_net_1 , N_149, 
        \crc_init_ff_RNO[13]_net_1 , N_144, \crc_unit_out[18] , 
        \crc_unit_out[13] , \buffer_ff_RNO[11]_net_1 , N_281, 
        \byte_ff_RNO[11]_net_1 , N_177, \crc_poly_ff_RNO[11]_net_1 , 
        N_209, \crc_out_ff[20]_net_1 , \buffer_ff[11]_net_1 , 
        \bus_reversed[11] , \crc_init_ff_3[8] , 
        \crc_poly_ff_RNO[24]_net_1 , N_222, \crc_init_ff_RNO[8]_net_1 , 
        N_139, \crc_poly_ff_RNO[8]_net_1 , N_206, 
        \crc_out_ff_RNO[5]_net_1 , N_243, \crc_out_ff_RNO[26]_net_1 , 
        N_264, \crc_unit_out[26] , \crc_unit_out[5] , N_244, 
        \crc_unit_out[6] , \crc_out_ff_RNO[6]_net_1 , 
        \crc_poly_ff_RNO[6]_net_1 , N_204, \crc_poly_ff_RNO[3]_net_1 , 
        N_201, \crc_idr_ff_RNO[6]_net_1 , N_236, 
        \crc_idr_ff_RNO[3]_net_1 , N_233, \crc_idr_ff_RNO[2]_net_1 , 
        N_232, \crc_poly_ff_RNO[2]_net_1 , N_200, \crc_init_mux[1] , 
        N_246, \crc_unit_out[8] , \crc_out_ff_RNO[8]_net_1 , N_274, 
        \bus_reversed[4] , \buffer_ff_RNO[4]_net_1 , N_262, 
        \crc_unit_out[24] , \crc_out_ff_RNO[24]_net_1 , 
        crc_poly_size_75_net_1, \crc_init_ff_3[7] , \crc_init_ff_3[0] , 
        \crc_init_ff_RNO[7]_net_1 , N_138, \crc_init_ff_RNO[0]_net_1 , 
        N_131, \crc_poly_ff_RNO[4]_net_1 , N_202, 
        \crc_out_ff_RNO[0]_net_1 , N_238, \crc_init_mux[23] , 
        \crc_init_mux[7] , \crc_unit_out[0] , N_157, 
        \crc_init_ff_3[26] , \crc_init_ff_RNO[26]_net_1 , N_252, 
        \crc_unit_out[14] , \crc_out_ff_RNO[14]_net_1 , 
        \crc_init_ff_3[14] , \crc_init_ff_3[30] , \crc_data_in0[6] , 
        \crc_data_in[6] , N_110, N_102, \byte_ff[30]_net_1 , 
        \byte_ff[14]_net_1 , \byte_ff[22]_net_1 , 
        \crc_out_ff_RNO[17]_net_1 , N_255, \crc_out_ff_RNO[30]_net_1 , 
        N_268, \buffer_ff_RNO[30]_net_1 , N_300, 
        \buffer_ff_RNO[22]_net_1 , N_292, \byte_ff_RNO[14]_net_1 , 
        N_180, \byte_ff_RNO[22]_net_1 , N_188, \byte_ff_RNO[30]_net_1 , 
        N_196, \crc_init_ff_RNO[14]_net_1 , N_145, 
        \crc_init_ff_RNO[30]_net_1 , N_161, \crc_init_mux[14] , 
        \crc_init_mux[6] , \crc_init_mux[30] , \buffer_ff[30]_net_1 , 
        \bus_reversed[30] , \buffer_ff[22]_net_1 , \bus_reversed[22] , 
        \crc_unit_out[30] , \crc_unit_out[17] , N_282, 
        \bus_reversed[12] , \buffer_ff_RNO[12]_net_1 , 
        \crc_init_ff_3[19] , \crc_out_ff_RNO[12]_net_1 , N_250, 
        \crc_out_ff_RNO[19]_net_1 , N_257, \crc_poly_ff_RNO[19]_net_1 , 
        N_217, \buffer_ff_RNO[20]_net_1 , N_290, 
        \byte_ff_RNO[20]_net_1 , N_186, \crc_init_ff_RNO[19]_net_1 , 
        N_150, \buffer_ff[20]_net_1 , \bus_reversed[20] , 
        \crc_unit_out[19] , \crc_unit_out[12] , N_249, 
        \crc_unit_out[11] , N_142, \crc_init_ff_3[11] , 
        \crc_init_ff_RNO[11]_net_1 , \crc_out_ff_RNO[11]_net_1 , N_210, 
        \crc_poly_ff_RNO[12]_net_1 , \crc_init_ff_3[12] , 
        \crc_init_ff_3[20] , \crc_out_ff_RNO[4]_net_1 , N_242, 
        \crc_out_ff_RNO[20]_net_1 , N_258, \crc_poly_ff_RNO[20]_net_1 , 
        N_218, \crc_init_ff_RNO[20]_net_1 , N_151, 
        \crc_init_ff_RNO[12]_net_1 , N_143, \crc_init_mux[20] , 
        \crc_unit_out[20] , \crc_unit_out[4] , GND, VCC;
    
    OR2A \crc_init_ff_RNO_1[20]  (.A(crc_init_en_0), .B(N_363), .Y(
        \crc_init_ff_3[20] ));
    NOR2B \crc_out_ff_RNO[21]  (.A(N_259), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[21]_net_1 ));
    MX2 \buffer_ff_RNO_0[14]  (.A(\buffer_ff[14]_net_1 ), .B(
        \bus_reversed[14] ), .S(buffer_en_0), .Y(N_284));
    OR2A \crc_init_ff_RNO_1[10]  (.A(crc_init_en_0), .B(N_353), .Y(
        \crc_init_ff_3[10] ));
    DFN1 \crc_init_ff[19]  (.D(\crc_init_ff_RNO[19]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[19]));
    DFN1 \crc_out_ff[13]  (.D(\crc_out_ff_RNO[13]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[13]_net_1 ));
    OR2A \byte_ff_RNO[20]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_186)
        , .Y(\byte_ff_RNO[20]_net_1 ));
    DFN1 \byte_ff[27]  (.D(\byte_ff_RNO[27]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[27]_net_1 ));
    DFN1 \byte_ff[24]  (.D(\byte_ff_RNO[24]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[24]_net_1 ));
    OR2A \crc_poly_ff_RNO[12]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_210), .Y(\crc_poly_ff_RNO[12]_net_1 ));
    OR2A \crc_init_ff_RNO_1[29]  (.A(crc_init_en), .B(N_335), .Y(
        \crc_init_ff_3[29] ));
    DFN1 \crc_init_ff[16]  (.D(\crc_init_ff_RNO[16]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[16]));
    DFN1 \buffer_ff[9]  (.D(\buffer_ff_RNO[9]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[9]_net_1 ));
    MX2 \crc_init_ff_RNO_0[13]  (.A(\crc_init_ff_3[13] ), .B(
        crc_init_out[13]), .S(un1_crc_init_en_1_0_net_1), .Y(N_144));
    OR2A \crc_init_ff_RNO_1[19]  (.A(crc_init_en_0), .B(N_362), .Y(
        \crc_init_ff_3[19] ));
    DFN1 \crc_idr_ff[6]  (.D(\crc_idr_ff_RNO[6]_net_1 ), .CLK(FAB_CLK), 
        .Q(crc_idr_out[6]));
    MX2 \crc_poly_ff_RNO_0[23]  (.A(crc_poly_out[23]), .B(N_366), .S(
        crc_poly_en_0), .Y(N_221));
    MX2 \bf_size_ff_RNO_0[0]  (.A(\bf_size_ff[0]_net_1 ), .B(
        \bf_size_ff_4[0] ), .S(un1_buffer_en_net_1), .Y(N_163));
    DFN1 \crc_init_ff[18]  (.D(\crc_init_ff_RNO[18]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[18]));
    DFN1 \crc_idr_ff[0]  (.D(\crc_idr_ff_RNO[0]_net_1 ), .CLK(FAB_CLK), 
        .Q(crc_idr_out[0]));
    MX2 \crc_init_ff_RNO_0[15]  (.A(\crc_init_ff_3[15] ), .B(
        crc_init_out[15]), .S(un1_crc_init_en_1_0_net_1), .Y(N_146));
    DFN1 \crc_out_ff[19]  (.D(\crc_out_ff_RNO[19]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[19]_net_1 ));
    MX2 \byte_ff_RNI15BP[14]  (.A(\byte_ff[30]_net_1 ), .B(
        \byte_ff[14]_net_1 ), .S(N_128), .Y(N_110));
    NOR2B \crc_poly_ff_RNO[21]  (.A(N_219), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[21]_net_1 ));
    NOR2B \crc_out_ff_RNO[4]  (.A(N_242), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[4]_net_1 ));
    DFN1 \crc_init_ff[13]  (.D(\crc_init_ff_RNO[13]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[13]));
    MX2 \crc_poly_ff_RNO_0[17]  (.A(crc_poly_out[17]), .B(N_360), .S(
        crc_poly_en_0), .Y(N_215));
    MX2 \byte_ff_RNO_0[29]  (.A(\byte_ff[29]_net_1 ), .B(
        \buffer_ff[29]_net_1 ), .S(byte_en), .Y(N_195));
    MX2 \buffer_ff_RNO_0[27]  (.A(\buffer_ff[27]_net_1 ), .B(
        \bus_reversed[27] ), .S(buffer_en), .Y(N_297));
    MX2 \byte_ff_RNIT3BA1[22]  (.A(\byte_ff[22]_net_1 ), .B(
        \crc_data_in0[6] ), .S(N_128), .Y(N_102));
    NOR2B \crc_poly_ff_RNO[29]  (.A(N_227), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[29]_net_1 ));
    NOR2B \crc_out_ff_RNO[6]  (.A(N_244), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[6]_net_1 ));
    DFN1 \crc_out_ff[15]  (.D(\crc_out_ff_RNO[15]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[15]_net_1 ));
    OR2A \crc_init_ff_RNO_1[2]  (.A(crc_init_en), .B(bus_wr_2), .Y(
        \crc_init_ff_3[2] ));
    NOR2B \crc_out_ff_RNO[19]  (.A(N_257), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[19]_net_1 ));
    MX2 \crc_out_ff_RNIR56K[8]  (.A(\crc_out_ff[23]_net_1 ), .B(
        \crc_out_ff[8]_net_1 ), .S(rev_out_type), .Y(crc_out[23]));
    MX2 \crc_init_ff_RNIS0EL[7]  (.A(crc_init_out[7]), .B(
        \crc_out_ff[7]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[7] ));
    DFN1 \crc_init_ff[3]  (.D(\crc_init_ff_RNO[3]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[3]));
    OR2A \byte_ff_RNO[6]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_172), 
        .Y(\byte_ff_RNO[6]_net_1 ));
    MX2 \byte_ff_RNO_0[11]  (.A(\byte_ff[11]_net_1 ), .B(
        \buffer_ff[11]_net_1 ), .S(byte_en_0), .Y(N_177));
    DFN1 \buffer_ff[0]  (.D(\buffer_ff_RNO[0]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[0]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[4]  (.A(crc_poly_out[4]), .B(N_347), .S(
        crc_poly_en), .Y(N_202));
    DFN1 \crc_poly_ff[12]  (.D(\crc_poly_ff_RNO[12]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[12]));
    MX2 \buffer_ff_RNO_0[5]  (.A(\buffer_ff[5]_net_1 ), .B(
        \bus_reversed[5] ), .S(buffer_en_0), .Y(N_275));
    MX2 \buffer_ff_RNO_0[16]  (.A(\buffer_ff[16]_net_1 ), .B(
        \bus_reversed[16] ), .S(buffer_en_0), .Y(N_286));
    MX2 \crc_init_ff_RNO_0[24]  (.A(\crc_init_ff_3[24] ), .B(
        crc_init_out[24]), .S(un1_crc_init_en_1_net_1), .Y(N_155));
    MX2 \buffer_ff_RNO_0[19]  (.A(\buffer_ff[19]_net_1 ), .B(
        \bus_reversed[19] ), .S(buffer_en), .Y(N_289));
    MX2 \crc_idr_ff_RNO_0[1]  (.A(crc_idr_out[1]), .B(bus_wr_1), .S(
        crc_idr_en), .Y(N_231));
    OR2A \buffer_ff_RNO[16]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_286), .Y(\buffer_ff_RNO[16]_net_1 ));
    NOR2B \bf_size_ff_RNO_1[0]  (.A(bus_size[0]), .B(buffer_en), .Y(
        \bf_size_ff_4[0] ));
    NOR2B \crc_poly_ff_RNO[30]  (.A(N_228), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[30]_net_1 ));
    OR2A \byte_ff_RNO[24]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_190)
        , .Y(\byte_ff_RNO[24]_net_1 ));
    MX2 \crc_out_ff_RNO_0[0]  (.A(\crc_unit_out[0] ), .B(
        \crc_out_ff[0]_net_1 ), .S(state_byte[4]), .Y(N_238));
    DFN1 \crc_poly_ff[20]  (.D(\crc_poly_ff_RNO[20]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[20]));
    OR2A \buffer_ff_RNO[15]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_285), .Y(\buffer_ff_RNO[15]_net_1 ));
    OR2A \buffer_ff_RNO[13]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_283), .Y(\buffer_ff_RNO[13]_net_1 ));
    MX2 \crc_init_ff_RNI22UR[28]  (.A(crc_init_out[28]), .B(
        \crc_out_ff[28]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[28] ));
    OR2A \bf_size_ff_RNO[1]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_164), .Y(\bf_size_ff_RNO[1]_net_1 ));
    OR2A \crc_poly_ff_RNO[22]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_220), .Y(\crc_poly_ff_RNO[22]_net_1 ));
    MX2 \crc_init_ff_RNIEIDL[0]  (.A(crc_init_out[0]), .B(
        \crc_out_ff[0]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[0] ));
    MX2 \buffer_ff_RNO_0[23]  (.A(\buffer_ff[23]_net_1 ), .B(
        \bus_reversed[23] ), .S(buffer_en), .Y(N_293));
    MX2 \byte_ff_RNO_0[18]  (.A(\byte_ff[18]_net_1 ), .B(
        \buffer_ff[18]_net_1 ), .S(byte_en), .Y(N_184));
    DFN1 \byte_ff[29]  (.D(\byte_ff_RNO[29]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[29]_net_1 ));
    OR2A \buffer_ff_RNO[12]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_282), .Y(\buffer_ff_RNO[12]_net_1 ));
    MX2 \crc_init_ff_RNIKODL[3]  (.A(crc_init_out[3]), .B(
        \crc_out_ff[3]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[3] ));
    OR2A \crc_init_ff_RNO[20]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_151), .Y(\crc_init_ff_RNO[20]_net_1 ));
    OR2A \crc_init_ff_RNO_1[1]  (.A(crc_init_en), .B(bus_wr_1), .Y(
        \crc_init_ff_3[1] ));
    MX2 \byte_ff_RNO_0[8]  (.A(\byte_ff[8]_net_1 ), .B(
        \buffer_ff[8]_net_1 ), .S(byte_en_0), .Y(N_174));
    OR2A \crc_init_ff_RNO_1[24]  (.A(crc_init_en_0), .B(N_367), .Y(
        \crc_init_ff_3[24] ));
    MX2 \crc_init_ff_RNO_0[30]  (.A(\crc_init_ff_3[30] ), .B(
        crc_init_out[30]), .S(un1_crc_init_en_1_net_1), .Y(N_161));
    DFN1 \byte_ff[16]  (.D(\byte_ff_RNO[16]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[16]_net_1 ));
    MX2 \byte_ff_RNINS9A1[17]  (.A(\byte_ff[17]_net_1 ), .B(
        \crc_data_in0[1] ), .S(N_128), .Y(N_97));
    DFN1 \crc_out_ff[0]  (.D(\crc_out_ff_RNO[0]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_out_ff[0]_net_1 ));
    OR2A \byte_ff_RNO[4]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_170), 
        .Y(\byte_ff_RNO[4]_net_1 ));
    DFN1 \buffer_ff[6]  (.D(\buffer_ff_RNO[6]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[6]_net_1 ));
    OR2A \crc_init_ff_RNO_1[14]  (.A(crc_init_en_0), .B(N_357), .Y(
        \crc_init_ff_3[14] ));
    MX2 \crc_init_ff_RNO_0[22]  (.A(\crc_init_ff_3[22] ), .B(
        crc_init_out[22]), .S(un1_crc_init_en_1_net_1), .Y(N_153));
    MX2 \crc_init_ff_RNIOU9Q[24]  (.A(crc_init_out[24]), .B(
        \crc_out_ff[24]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[24] ));
    DFN1 \buffer_ff[19]  (.D(\buffer_ff_RNO[19]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[19]_net_1 ));
    OR2A \byte_ff_RNO[13]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_179)
        , .Y(\byte_ff_RNO[13]_net_1 ));
    DFN1 \byte_ff[2]  (.D(\byte_ff_RNO[2]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[2]_net_1 ));
    OR2A \crc_init_ff_RNO[23]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_154), .Y(\crc_init_ff_RNO[23]_net_1 ));
    NOR2B \crc_out_ff_RNO[28]  (.A(N_266), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[28]_net_1 ));
    MX2 \byte_ff_RNIIAIL[0]  (.A(\byte_ff[0]_net_1 ), .B(
        \buffer_ff[0]_net_1 ), .S(bypass_byte0), .Y(\crc_data_in0[0] ));
    MX2 \byte_ff_RNO_0[22]  (.A(\byte_ff[22]_net_1 ), .B(
        \buffer_ff[22]_net_1 ), .S(byte_en), .Y(N_188));
    MX2 \crc_out_ff_RNO_0[9]  (.A(\crc_unit_out[9] ), .B(
        \crc_out_ff[9]_net_1 ), .S(state_byte[4]), .Y(N_247));
    OR2A \crc_init_ff_RNO_1[4]  (.A(crc_init_en), .B(N_347), .Y(
        \crc_init_ff_3[4] ));
    OR2A \crc_init_ff_RNO[26]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_157), .Y(\crc_init_ff_RNO[26]_net_1 ));
    MX2 \byte_ff_RNO_0[9]  (.A(\byte_ff[9]_net_1 ), .B(
        \buffer_ff[9]_net_1 ), .S(byte_en_0), .Y(N_175));
    MX2 \byte_ff_RNO_0[27]  (.A(\byte_ff[27]_net_1 ), .B(
        \buffer_ff[27]_net_1 ), .S(byte_en), .Y(N_193));
    OR2A \byte_ff_RNO[18]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_184)
        , .Y(\byte_ff_RNO[18]_net_1 ));
    MX2 \buffer_ff_RNO_0[12]  (.A(\buffer_ff[12]_net_1 ), .B(
        \bus_reversed[12] ), .S(buffer_en_0), .Y(N_282));
    DFN1 \size_ff[1]  (.D(\size_ff_RNO[1]_net_1 ), .CLK(FAB_CLK), .Q(
        \size_ff[1]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[2]  (.A(crc_poly_out[2]), .B(bus_wr_2), .S(
        crc_poly_en), .Y(N_200));
    MX2 \crc_poly_ff_RNO_0[21]  (.A(crc_poly_out[21]), .B(N_364), .S(
        crc_poly_en_0), .Y(N_219));
    NOR2B \crc_out_ff_RNO[17]  (.A(N_255), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[17]_net_1 ));
    OR2A \crc_init_ff_RNO_1[30]  (.A(crc_init_en), .B(N_336), .Y(
        \crc_init_ff_3[30] ));
    OR2A \crc_init_ff_RNO_1[22]  (.A(crc_init_en_0), .B(N_365), .Y(
        \crc_init_ff_3[22] ));
    OR2A \crc_init_ff_RNO[17]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_148), .Y(\crc_init_ff_RNO[17]_net_1 ));
    MX2 \crc_out_ff_RNIIT6K[0]  (.A(\crc_out_ff[31]_net_1 ), .B(
        \crc_out_ff[0]_net_1 ), .S(rev_out_type), .Y(crc_out[31]));
    DFN1 \byte_ff[20]  (.D(\byte_ff_RNO[20]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[20]_net_1 ));
    MX2 \crc_out_ff_RNO_0[5]  (.A(\crc_unit_out[5] ), .B(
        \crc_out_ff[5]_net_1 ), .S(state_byte[4]), .Y(N_243));
    DFN1 \crc_init_ff[25]  (.D(\crc_init_ff_RNO[25]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[25]));
    DFN1 \byte_ff[17]  (.D(\byte_ff_RNO[17]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[17]_net_1 ));
    DFN1 \byte_ff[14]  (.D(\byte_ff_RNO[14]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[14]_net_1 ));
    NOR2B \crc_out_ff_RNO[12]  (.A(N_250), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[12]_net_1 ));
    OR2A \crc_init_ff_RNO_1[12]  (.A(crc_init_en_0), .B(N_355), .Y(
        \crc_init_ff_3[12] ));
    MX2 \crc_poly_ff_RNO_0[7]  (.A(crc_poly_out[7]), .B(N_350), .S(
        crc_poly_en), .Y(N_205));
    MX2 \byte_ff_RNITTPJ2[11]  (.A(N_107), .B(N_99), .S(N_294_0), .Y(
        \crc_data_in[3] ));
    DFN1 \buffer_ff[7]  (.D(\buffer_ff_RNO[7]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[7]_net_1 ));
    OR2A \byte_ff_RNO[0]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_166), 
        .Y(\byte_ff_RNO[0]_net_1 ));
    OR2A \crc_init_ff_RNO[2]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_133), .Y(\crc_init_ff_RNO[2]_net_1 ));
    OR2A \buffer_ff_RNO[29]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_299), .Y(\buffer_ff_RNO[29]_net_1 ));
    OR2A \crc_poly_ff_RNO[0]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_198), .Y(\crc_poly_ff_RNO[0]_net_1 ));
    DFN1 \crc_poly_ff[19]  (.D(\crc_poly_ff_RNO[19]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[19]));
    MX2 \crc_poly_ff_RNO_0[15]  (.A(crc_poly_out[15]), .B(N_358), .S(
        crc_poly_en_0), .Y(N_213));
    OR2A \buffer_ff_RNO[2]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_272), .Y(\buffer_ff_RNO[2]_net_1 ));
    MX2 \crc_init_ff_RNIS2AQ[26]  (.A(crc_init_out[26]), .B(
        \crc_out_ff[26]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[26] ));
    MX2 \byte_ff_RNI0PIL[7]  (.A(\byte_ff[7]_net_1 ), .B(
        \buffer_ff[7]_net_1 ), .S(bypass_byte0), .Y(\crc_data_in0[7] ));
    OR2A \buffer_ff_RNO[20]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_290), .Y(\buffer_ff_RNO[20]_net_1 ));
    DFN1 \crc_out_ff[20]  (.D(\crc_out_ff_RNO[20]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[20]_net_1 ));
    MX2 \buffer_ff_RNO_0[20]  (.A(\buffer_ff[20]_net_1 ), .B(
        \bus_reversed[20] ), .S(buffer_en), .Y(N_290));
    DFN1 \crc_out_ff[21]  (.D(\crc_out_ff_RNO[21]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[21]_net_1 ));
    MX2 \crc_init_ff_RNI44UR[29]  (.A(crc_init_out[29]), .B(
        \crc_out_ff[29]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[29] ));
    DFN1 \crc_out_ff[3]  (.D(\crc_out_ff_RNO[3]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_out_ff[3]_net_1 ));
    DFN1 \byte_ff[5]  (.D(\byte_ff_RNO[5]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[5]_net_1 ));
    MX2 \crc_init_ff_RNIU2EL[8]  (.A(crc_init_out[8]), .B(
        \crc_out_ff[8]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[8] ));
    MX2 \crc_out_ff_RNI2RHQ[11]  (.A(\crc_out_ff[20]_net_1 ), .B(
        \crc_out_ff[11]_net_1 ), .S(rev_out_type), .Y(crc_out[20]));
    NOR2B \crc_poly_ff_RNO[13]  (.A(N_211), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[13]_net_1 ));
    OR2A \buffer_ff_RNO[27]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_297), .Y(\buffer_ff_RNO[27]_net_1 ));
    DFN1 \crc_out_ff[22]  (.D(\crc_out_ff_RNO[22]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[22]_net_1 ));
    MX2 \byte_ff_RNO_0[19]  (.A(\byte_ff[19]_net_1 ), .B(
        \buffer_ff[19]_net_1 ), .S(byte_en), .Y(N_185));
    OR2A \crc_init_ff_RNO[9]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_140), .Y(\crc_init_ff_RNO[9]_net_1 ));
    NOR2B \crc_out_ff_RNO[25]  (.A(N_263), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[25]_net_1 ));
    OR2A \crc_init_ff_RNO[31]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_162), .Y(\crc_init_ff_RNO[31]_net_1 ));
    DFN1 \crc_out_ff[26]  (.D(\crc_out_ff_RNO[26]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[26]_net_1 ));
    MX2 \crc_out_ff_RNO_0[24]  (.A(\crc_unit_out[24] ), .B(
        \crc_out_ff[24]_net_1 ), .S(state_byte_0[4]), .Y(N_262));
    DFN1 \buffer_ff[12]  (.D(\buffer_ff_RNO[12]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[12]_net_1 ));
    NOR2A crc_poly_size_76_1 (.A(crc_poly_size[0]), .B(
        crc_poly_size[1]), .Y(crc_poly_size_76_1_net_1));
    OR2A \crc_poly_ff_RNO[16]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_214), .Y(\crc_poly_ff_RNO[16]_net_1 ));
    MX2 \crc_out_ff_RNO_0[16]  (.A(\crc_unit_out[16] ), .B(
        \crc_out_ff[16]_net_1 ), .S(state_byte_0[4]), .Y(N_254));
    MX2 \crc_init_ff_RNIKO7Q[13]  (.A(crc_init_out[13]), .B(
        \crc_out_ff[13]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[13] ));
    MX2 \crc_init_ff_RNO_0[21]  (.A(\crc_init_ff_3[21] ), .B(
        crc_init_out[21]), .S(un1_crc_init_en_1_net_1), .Y(N_152));
    MX2 \crc_out_ff_RNO_0[7]  (.A(\crc_unit_out[7] ), .B(
        \crc_out_ff[7]_net_1 ), .S(state_byte[4]), .Y(N_245));
    NOR2B \crc_idr_ff_RNO[7]  (.A(N_237), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_idr_ff_RNO[7]_net_1 ));
    OR2A \crc_init_ff_RNO[24]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_155), .Y(\crc_init_ff_RNO[24]_net_1 ));
    DFN1 \crc_out_ff[17]  (.D(\crc_out_ff_RNO[17]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[17]_net_1 ));
    DFN1 \buffer_ff[29]  (.D(\buffer_ff_RNO[29]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[29]_net_1 ));
    DFN1 \byte_ff[4]  (.D(\byte_ff_RNO[4]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[4]_net_1 ));
    DFN1 \byte_ff[7]  (.D(\byte_ff_RNO[7]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[7]_net_1 ));
    DFN1 \byte_ff[19]  (.D(\byte_ff_RNO[19]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[19]_net_1 ));
    MX2 \crc_out_ff_RNO_0[15]  (.A(\crc_unit_out[15] ), .B(
        \crc_out_ff[15]_net_1 ), .S(state_byte_0[4]), .Y(N_253));
    DFN1 \byte_ff[6]  (.D(\byte_ff_RNO[6]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[6]_net_1 ));
    MX2 \crc_out_ff_RNIB3HQ[12]  (.A(\crc_out_ff[19]_net_1 ), .B(
        \crc_out_ff[12]_net_1 ), .S(rev_out_type), .Y(crc_out[19]));
    DFN1 \crc_out_ff[28]  (.D(\crc_out_ff_RNO[28]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[28]_net_1 ));
    OR2A \crc_init_ff_RNO[28]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_159), .Y(\crc_init_ff_RNO[28]_net_1 ));
    DFN1 \crc_out_ff[2]  (.D(\crc_out_ff_RNO[2]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_out_ff[2]_net_1 ));
    OR2A \byte_ff_RNO[23]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_189)
        , .Y(\byte_ff_RNO[23]_net_1 ));
    MX2 \buffer_ff_RNO_0[21]  (.A(\buffer_ff[21]_net_1 ), .B(
        \bus_reversed[21] ), .S(buffer_en), .Y(N_291));
    MX2 \crc_init_ff_RNO_0[10]  (.A(\crc_init_ff_3[10] ), .B(
        crc_init_out[10]), .S(un1_crc_init_en_1_0_net_1), .Y(N_141));
    MX2 \byte_ff_RNI7KAH2[8]  (.A(N_104), .B(N_96), .S(N_294_0), .Y(
        \crc_data_in[0] ));
    MX2 \buffer_ff_RNO_0[8]  (.A(\buffer_ff[8]_net_1 ), .B(
        \bus_reversed[8] ), .S(buffer_en_0), .Y(N_278));
    MX2 \byte_ff_RNO_0[7]  (.A(\byte_ff[7]_net_1 ), .B(
        \buffer_ff[7]_net_1 ), .S(byte_en_0), .Y(N_173));
    MX2 \crc_out_ff_RNIR56K[7]  (.A(\crc_out_ff[24]_net_1 ), .B(
        \crc_out_ff[7]_net_1 ), .S(rev_out_type), .Y(crc_out[24]));
    DFN1 \crc_poly_ff[0]  (.D(\crc_poly_ff_RNO[0]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[0]));
    DFN1 \crc_poly_ff[5]  (.D(\crc_poly_ff_RNO[5]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[5]));
    OR2A \byte_ff_RNO[2]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_168), 
        .Y(\byte_ff_RNO[2]_net_1 ));
    OR2A \byte_ff_RNO[28]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_194)
        , .Y(\byte_ff_RNO[28]_net_1 ));
    DFN1 \crc_poly_ff[25]  (.D(\crc_poly_ff_RNO[25]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[25]));
    MX2 \crc_out_ff_RNIR56K[9]  (.A(\crc_out_ff[22]_net_1 ), .B(
        \crc_out_ff[9]_net_1 ), .S(rev_out_type), .Y(crc_out[22]));
    MX2 \byte_ff_RNIP8RM[9]  (.A(\byte_ff[25]_net_1 ), .B(
        \byte_ff[9]_net_1 ), .S(N_128), .Y(N_105));
    MX2 \crc_poly_ff_RNO_0[8]  (.A(crc_poly_out[8]), .B(N_351), .S(
        crc_poly_en), .Y(N_206));
    DFN1 \buffer_ff[11]  (.D(\buffer_ff_RNO[11]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[11]_net_1 ));
    DFN1 \byte_ff[23]  (.D(\byte_ff_RNO[23]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[23]_net_1 ));
    OR2A \buffer_ff_RNO[30]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_300), .Y(\buffer_ff_RNO[30]_net_1 ));
    DFN1 \buffer_ff[17]  (.D(\buffer_ff_RNO[17]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[17]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[18]  (.A(crc_poly_out[18]), .B(N_361), .S(
        crc_poly_en_0), .Y(N_216));
    OR2A \crc_poly_ff_RNO[23]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_221), .Y(\crc_poly_ff_RNO[23]_net_1 ));
    OR2A \crc_init_ff_RNO_1[21]  (.A(crc_init_en_0), .B(N_364), .Y(
        \crc_init_ff_3[21] ));
    OR2A \crc_init_ff_RNO[22]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_153), .Y(\crc_init_ff_RNO[22]_net_1 ));
    MX2 \crc_init_ff_RNO_0[19]  (.A(\crc_init_ff_3[19] ), .B(
        crc_init_out[19]), .S(un1_crc_init_en_1_net_1), .Y(N_150));
    DFN1 \bf_size_ff[0]  (.D(\bf_size_ff_RNO[0]_net_1 ), .CLK(FAB_CLK), 
        .Q(\bf_size_ff[0]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1 \crc_poly_ff[3]  (.D(\crc_poly_ff_RNO[3]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[3]));
    MX2 \crc_out_ff_RNO_0[6]  (.A(\crc_unit_out[6] ), .B(
        \crc_out_ff[6]_net_1 ), .S(state_byte[4]), .Y(N_244));
    MX2 \crc_out_ff_RNO_0[23]  (.A(\crc_unit_out[23] ), .B(
        \crc_out_ff[23]_net_1 ), .S(state_byte_0[4]), .Y(N_261));
    NOR2B \crc_out_ff_RNO[31]  (.A(N_269), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[31]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[10]  (.A(crc_poly_out[10]), .B(N_353), .S(
        crc_poly_en_0), .Y(N_208));
    OR2A \crc_init_ff_RNO_1[11]  (.A(crc_init_en_0), .B(N_354), .Y(
        \crc_init_ff_3[11] ));
    DFN1 \crc_poly_ff[21]  (.D(\crc_poly_ff_RNO[21]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[21]));
    DFN1 \crc_poly_ff[10]  (.D(\crc_poly_ff_RNO[10]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[10]));
    DFN1 \crc_out_ff[6]  (.D(\crc_out_ff_RNO[6]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_out_ff[6]_net_1 ));
    MX2 \crc_init_ff_RNO_0[9]  (.A(\crc_init_ff_3[9] ), .B(
        crc_init_out[9]), .S(un1_crc_init_en_1_0_net_1), .Y(N_140));
    OR2A \crc_poly_ff_RNO[26]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_224), .Y(\crc_poly_ff_RNO[26]_net_1 ));
    MX2 \crc_init_ff_RNIQ0AQ[25]  (.A(crc_init_out[25]), .B(
        \crc_out_ff[25]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[25] ));
    DFN1 \byte_ff[25]  (.D(\byte_ff_RNO[25]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[25]_net_1 ));
    MX2 \buffer_ff_RNO_0[24]  (.A(\buffer_ff[24]_net_1 ), .B(
        \bus_reversed[24] ), .S(buffer_en), .Y(N_294));
    DFN1 \crc_out_ff[23]  (.D(\crc_out_ff_RNO[23]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[23]_net_1 ));
    MX2 \byte_ff_RNO_0[12]  (.A(\byte_ff[12]_net_1 ), .B(
        \buffer_ff[12]_net_1 ), .S(byte_en_0), .Y(N_178));
    MX2 \byte_ff_RNI47AP[11]  (.A(\byte_ff[27]_net_1 ), .B(
        \byte_ff[11]_net_1 ), .S(N_128), .Y(N_107));
    MX2 \byte_ff_RNO_0[17]  (.A(\byte_ff[17]_net_1 ), .B(
        \buffer_ff[17]_net_1 ), .S(byte_en), .Y(N_183));
    MX2 \crc_out_ff_RNI92IL[12]  (.A(\crc_out_ff[12]_net_1 ), .B(
        \crc_out_ff[19]_net_1 ), .S(rev_out_type_0), .Y(crc_out[12]));
    MX2 \crc_out_ff_RNO_0[31]  (.A(\crc_unit_out[31] ), .B(
        \crc_out_ff[31]_net_1 ), .S(state_byte[4]), .Y(N_269));
    OR2A \byte_ff_RNO[3]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_169), 
        .Y(\byte_ff_RNO[3]_net_1 ));
    MX2 \buffer_ff_RNO_0[1]  (.A(\buffer_ff[1]_net_1 ), .B(
        \bus_reversed[1] ), .S(buffer_en_0), .Y(N_271));
    MX2 \byte_ff_RNO_0[23]  (.A(\byte_ff[23]_net_1 ), .B(
        \buffer_ff[23]_net_1 ), .S(byte_en), .Y(N_189));
    DFN1 \crc_poly_ff[7]  (.D(\crc_poly_ff_RNO[7]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[7]));
    OR2A \buffer_ff_RNO[5]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_275), .Y(\buffer_ff_RNO[5]_net_1 ));
    OR2A \crc_poly_ff_RNO[5]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_203), .Y(\crc_poly_ff_RNO[5]_net_1 ));
    OR2A \crc_init_ff_RNO[8]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_139), .Y(\crc_init_ff_RNO[8]_net_1 ));
    NOR2B \crc_out_ff_RNO[29]  (.A(N_267), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[29]_net_1 ));
    DFN1 \byte_ff[10]  (.D(\byte_ff_RNO[10]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[10]_net_1 ));
    OR2A \byte_ff_RNO[16]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_182)
        , .Y(\byte_ff_RNO[16]_net_1 ));
    DFN1 \crc_out_ff[5]  (.D(\crc_out_ff_RNO[5]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_out_ff[5]_net_1 ));
    NOR2B \crc_poly_ff_RNO[9]  (.A(N_207), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[9]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[19]  (.A(crc_poly_out[19]), .B(N_362), .S(
        crc_poly_en_0), .Y(N_217));
    OR2A \crc_init_ff_RNO[19]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_150), .Y(\crc_init_ff_RNO[19]_net_1 ));
    NOR2B \crc_out_ff_RNO[14]  (.A(N_252), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[14]_net_1 ));
    DFN1 \crc_init_ff[20]  (.D(\crc_init_ff_RNO[20]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[20]));
    OR2A \crc_init_ff_RNO[30]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_161), .Y(\crc_init_ff_RNO[30]_net_1 ));
    DFN1 \crc_poly_ff[27]  (.D(\crc_poly_ff_RNO[27]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[27]));
    DFN1 \crc_out_ff[29]  (.D(\crc_out_ff_RNO[29]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[29]_net_1 ));
    NOR2A crc_poly_size_75 (.A(crc_poly_size[1]), .B(crc_poly_size[0]), 
        .Y(crc_poly_size_75_net_1));
    DFN1 \crc_out_ff[25]  (.D(\crc_out_ff_RNO[25]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[25]_net_1 ));
    MX2 \byte_ff_RNIKCIL[1]  (.A(\byte_ff[1]_net_1 ), .B(
        \buffer_ff[1]_net_1 ), .S(bypass_byte0), .Y(\crc_data_in0[1] ));
    DFN1 \buffer_ff[22]  (.D(\buffer_ff_RNO[22]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[22]_net_1 ));
    OR2A \byte_ff_RNO[11]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_177)
        , .Y(\byte_ff_RNO[11]_net_1 ));
    MX2 \crc_out_ff_RNIIT6K[1]  (.A(\crc_out_ff[30]_net_1 ), .B(
        \crc_out_ff[1]_net_1 ), .S(rev_out_type), .Y(crc_out[30]));
    OR2A \buffer_ff_RNO[3]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_273), .Y(\buffer_ff_RNO[3]_net_1 ));
    MX2 \buffer_ff_RNO_0[26]  (.A(\buffer_ff[26]_net_1 ), .B(
        \bus_reversed[26] ), .S(buffer_en), .Y(N_296));
    MX2 \buffer_ff_RNO_0[29]  (.A(\buffer_ff[29]_net_1 ), .B(
        \bus_reversed[29] ), .S(buffer_en), .Y(N_299));
    MX2 \size_ff_RNO_0[1]  (.A(\size_ff[1]_net_1 ), .B(
        \bf_size_ff[1]_net_1 ), .S(byte_en_0), .Y(N_130));
    MX2 \size_ff_RNI5F3P[0]  (.A(\size_ff[0]_net_1 ), .B(
        \bf_size_ff[0]_net_1 ), .S(N_118_1), .Y(size_in[0]));
    DFN1 \crc_poly_ff[28]  (.D(\crc_poly_ff_RNO[28]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[28]));
    MX2 \crc_init_ff_RNO_0[14]  (.A(\crc_init_ff_3[14] ), .B(
        crc_init_out[14]), .S(un1_crc_init_en_1_0_net_1), .Y(N_145));
    OR2A \buffer_ff_RNO[28]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_298), .Y(\buffer_ff_RNO[28]_net_1 ));
    MX2 \crc_out_ff_RNIP47F[3]  (.A(\crc_out_ff[3]_net_1 ), .B(
        \crc_out_ff[28]_net_1 ), .S(rev_out_type_0), .Y(crc_out[3]));
    NOR2B \crc_poly_ff_RNO[14]  (.A(N_212), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[14]_net_1 ));
    DFN1 \crc_init_ff[6]  (.D(\crc_init_ff_RNO[6]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[6]));
    NOR2B \crc_idr_ff_RNO[2]  (.A(N_232), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_idr_ff_RNO[2]_net_1 ));
    DFN1 \crc_poly_ff[23]  (.D(\crc_poly_ff_RNO[23]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[23]));
    MX2 \buffer_ff_RNO_0[9]  (.A(\buffer_ff[9]_net_1 ), .B(
        \bus_reversed[9] ), .S(buffer_en_0), .Y(N_279));
    MX2 \crc_poly_ff_RNO_0[16]  (.A(crc_poly_out[16]), .B(bus_wr_16), 
        .S(crc_poly_en_0), .Y(N_214));
    MX2 \crc_out_ff_RNO_0[11]  (.A(\crc_unit_out[11] ), .B(
        \crc_out_ff[11]_net_1 ), .S(state_byte_0[4]), .Y(N_249));
    MX2 \crc_init_ff_RNIQU7Q[16]  (.A(crc_init_out[16]), .B(
        \crc_out_ff[16]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[16] ));
    MX2 \crc_idr_ff_RNO_0[4]  (.A(crc_idr_out[4]), .B(N_347), .S(
        crc_idr_en), .Y(N_234));
    OR2A \byte_ff_RNO[12]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_178)
        , .Y(\byte_ff_RNO[12]_net_1 ));
    NOR2B \crc_idr_ff_RNO[3]  (.A(N_233), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_idr_ff_RNO[3]_net_1 ));
    MX2 \crc_init_ff_RNO_0[31]  (.A(\crc_init_ff_3[31] ), .B(
        crc_init_out[31]), .S(un1_crc_init_en_1_net_1), .Y(N_162));
    DFN1 \buffer_ff[21]  (.D(\buffer_ff_RNO[21]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[21]_net_1 ));
    MX2 \byte_ff_RNIN6RM[8]  (.A(\byte_ff[24]_net_1 ), .B(
        \byte_ff[8]_net_1 ), .S(N_128), .Y(N_104));
    MX2 \crc_init_ff_RNIOSDL[5]  (.A(crc_init_out[5]), .B(
        \crc_out_ff[5]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[5] ));
    DFN1 \buffer_ff[27]  (.D(\buffer_ff_RNO[27]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[27]_net_1 ));
    MX2 \byte_ff_RNO_0[4]  (.A(\byte_ff[4]_net_1 ), .B(
        \buffer_ff[4]_net_1 ), .S(byte_en_0), .Y(N_170));
    MX2 \buffer_ff_RNO_0[30]  (.A(\buffer_ff[30]_net_1 ), .B(
        \bus_reversed[30] ), .S(buffer_en), .Y(N_300));
    MX2 \crc_out_ff_RNO_0[27]  (.A(\crc_unit_out[27] ), .B(
        \crc_out_ff[27]_net_1 ), .S(state_byte[4]), .Y(N_265));
    MX2 \crc_init_ff_RNIGKDL[1]  (.A(crc_init_out[1]), .B(
        \crc_out_ff[1]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[1] ));
    NOR2B \crc_out_ff_RNO[27]  (.A(N_265), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[27]_net_1 ));
    MX2 \crc_out_ff_RNIR56K[6]  (.A(\crc_out_ff[25]_net_1 ), .B(
        \crc_out_ff[6]_net_1 ), .S(rev_out_type), .Y(crc_out[25]));
    MX2 \crc_poly_ff_RNO_0[12]  (.A(crc_poly_out[12]), .B(N_355), .S(
        crc_poly_en_0), .Y(N_210));
    MX2 \crc_init_ff_RNIKQ9Q[22]  (.A(crc_init_out[22]), .B(
        \crc_out_ff[22]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[22] ));
    DFN1 \crc_init_ff[22]  (.D(\crc_init_ff_RNO[22]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[22]));
    MX2 \buffer_ff_RNO_0[4]  (.A(\buffer_ff[4]_net_1 ), .B(
        \bus_reversed[4] ), .S(buffer_en_0), .Y(N_274));
    MX2 \byte_ff_RNO_0[20]  (.A(\byte_ff[20]_net_1 ), .B(
        \buffer_ff[20]_net_1 ), .S(byte_en), .Y(N_186));
    MX2 \crc_poly_ff_RNO_0[6]  (.A(crc_poly_out[6]), .B(N_349), .S(
        crc_poly_en), .Y(N_204));
    MX2 \byte_ff_RNIUMIL[6]  (.A(\byte_ff[6]_net_1 ), .B(
        \buffer_ff[6]_net_1 ), .S(bypass_byte0), .Y(\crc_data_in0[6] ));
    MX2 \crc_out_ff_RNO_0[22]  (.A(\crc_unit_out[22] ), .B(
        \crc_out_ff[22]_net_1 ), .S(state_byte_0[4]), .Y(N_260));
    OR2A \crc_init_ff_RNO[11]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_142), .Y(\crc_init_ff_RNO[11]_net_1 ));
    MX2 \crc_init_ff_RNO_0[12]  (.A(\crc_init_ff_3[12] ), .B(
        crc_init_out[12]), .S(un1_crc_init_en_1_0_net_1), .Y(N_143));
    MX2 \crc_out_ff_RNO_0[8]  (.A(\crc_unit_out[8] ), .B(
        \crc_out_ff[8]_net_1 ), .S(state_byte[4]), .Y(N_246));
    MX2 \crc_init_ff_RNIKLVR[30]  (.A(crc_init_out[30]), .B(
        \crc_out_ff[30]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[30] ));
    DFN1 \byte_ff[13]  (.D(\byte_ff_RNO[13]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[13]_net_1 ));
    NOR2B \crc_out_ff_RNO[22]  (.A(N_260), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[22]_net_1 ));
    OA1A crc_init_sel_ff_RNIEJTVA (.A(state_byte_i[0]), .B(
        crc_init_sel_ff_net_1), .C(N_56), .Y(N_165));
    OR2A \byte_ff_RNO[19]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_185)
        , .Y(\byte_ff_RNO[19]_net_1 ));
    OR2A \buffer_ff_RNO[9]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_279), .Y(\buffer_ff_RNO[9]_net_1 ));
    DFN1 \crc_init_ff[21]  (.D(\crc_init_ff_RNO[21]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[21]));
    OR2A \crc_init_ff_RNO_1[31]  (.A(crc_init_en), .B(N_337), .Y(
        \crc_init_ff_3[31] ));
    MX2 \buffer_ff_RNO_0[22]  (.A(\buffer_ff[22]_net_1 ), .B(
        \bus_reversed[22] ), .S(buffer_en), .Y(N_292));
    NOR2B \crc_poly_ff_RNO[24]  (.A(N_222), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[24]_net_1 ));
    OR2A \byte_ff_RNO[26]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_192)
        , .Y(\byte_ff_RNO[26]_net_1 ));
    DFN1 \bf_size_ff[1]  (.D(\bf_size_ff_RNO[1]_net_1 ), .CLK(FAB_CLK), 
        .Q(\bf_size_ff[1]_net_1 ));
    MX2 \crc_out_ff_RNO_0[19]  (.A(\crc_unit_out[19] ), .B(
        \crc_out_ff[19]_net_1 ), .S(state_byte_0[4]), .Y(N_257));
    MX2 \crc_out_ff_RNO_0[18]  (.A(\crc_unit_out[18] ), .B(
        \crc_out_ff[18]_net_1 ), .S(state_byte_0[4]), .Y(N_256));
    NOR2B \crc_poly_ff_RNO[31]  (.A(N_229), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[31]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[30]  (.A(crc_poly_out[30]), .B(N_336), .S(
        crc_poly_en), .Y(N_228));
    MX2 \crc_poly_ff_RNO_0[14]  (.A(crc_poly_out[14]), .B(N_357), .S(
        crc_poly_en_0), .Y(N_212));
    OR2A \crc_init_ff_RNO_1[3]  (.A(crc_init_en), .B(bus_wr_3), .Y(
        \crc_init_ff_3[3] ));
    MX2 \crc_init_ff_RNO_0[0]  (.A(\crc_init_ff_3[0] ), .B(
        crc_init_out[0]), .S(un1_crc_init_en_1_0_net_1), .Y(N_131));
    DFN1 \byte_ff[15]  (.D(\byte_ff_RNO[15]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[15]_net_1 ));
    MX2 \crc_out_ff_RNI0QIL[10]  (.A(\crc_out_ff[10]_net_1 ), .B(
        \crc_out_ff[21]_net_1 ), .S(rev_out_type_0), .Y(crc_out[10]));
    NOR2B crc_poly_size_74 (.A(crc_poly_size[1]), .B(crc_poly_size[0]), 
        .Y(crc_poly_size_74_net_1));
    DFN1 \crc_init_ff[27]  (.D(\crc_init_ff_RNO[27]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[27]));
    MX2 \buffer_ff_RNO_0[31]  (.A(\buffer_ff[31]_net_1 ), .B(
        \bus_reversed[31] ), .S(buffer_en), .Y(N_301));
    NOR2B \crc_out_ff_RNO[13]  (.A(N_251), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[13]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[27]  (.A(crc_poly_out[27]), .B(N_333), .S(
        crc_poly_en), .Y(N_225));
    OR2A \buffer_ff_RNO[19]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_289), .Y(\buffer_ff_RNO[19]_net_1 ));
    NOR2B \crc_out_ff_RNO[8]  (.A(N_246), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[8]_net_1 ));
    MX2 \byte_ff_RNO_0[1]  (.A(\byte_ff[1]_net_1 ), .B(
        \buffer_ff[1]_net_1 ), .S(byte_en_0), .Y(N_167));
    MX2 \crc_out_ff_RNIGS7F[1]  (.A(\crc_out_ff[1]_net_1 ), .B(
        \crc_out_ff[30]_net_1 ), .S(rev_out_type_0), .Y(crc_out[1]));
    MX2 \byte_ff_RNO_0[31]  (.A(\byte_ff[31]_net_1 ), .B(
        \buffer_ff[31]_net_1 ), .S(byte_en), .Y(N_197));
    OR2A \buffer_ff_RNO[10]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_280), .Y(\buffer_ff_RNO[10]_net_1 ));
    MX2 \byte_ff_RNO_0[13]  (.A(\byte_ff[13]_net_1 ), .B(
        \buffer_ff[13]_net_1 ), .S(byte_en_0), .Y(N_179));
    MX2 \byte_ff_RNIKP9A1[16]  (.A(\byte_ff[16]_net_1 ), .B(
        \crc_data_in0[0] ), .S(N_128), .Y(N_96));
    MX2 \crc_poly_ff_RNO_0[1]  (.A(crc_poly_out[1]), .B(bus_wr_1), .S(
        crc_poly_en), .Y(N_199));
    OR2A \byte_ff_RNO[21]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_187)
        , .Y(\byte_ff_RNO[21]_net_1 ));
    MX2 \byte_ff_RNO_0[25]  (.A(\byte_ff[25]_net_1 ), .B(
        \buffer_ff[25]_net_1 ), .S(byte_en), .Y(N_191));
    DFN1 \byte_ff[21]  (.D(\byte_ff_RNO[21]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[21]_net_1 ));
    MX2 \byte_ff_RNO_0[26]  (.A(\byte_ff[26]_net_1 ), .B(
        \buffer_ff[26]_net_1 ), .S(byte_en), .Y(N_192));
    OR2A \size_ff_RNO[1]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_130), 
        .Y(\size_ff_RNO[1]_net_1 ));
    DFN1 \crc_poly_ff[15]  (.D(\crc_poly_ff_RNO[15]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[15]));
    NOR2B \crc_out_ff_RNO[3]  (.A(N_241), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[3]_net_1 ));
    MX2 \byte_ff_RNIOOPJ2[10]  (.A(N_106), .B(N_98), .S(N_294_0), .Y(
        \crc_data_in[2] ));
    MX2 \crc_init_ff_RNO_0[26]  (.A(\crc_init_ff_3[26] ), .B(
        crc_init_out[26]), .S(un1_crc_init_en_1_net_1), .Y(N_157));
    MX2 \byte_ff_RNO_0[5]  (.A(\byte_ff[5]_net_1 ), .B(
        \buffer_ff[5]_net_1 ), .S(byte_en_0), .Y(N_171));
    DFN1 \buffer_ff[5]  (.D(\buffer_ff_RNO[5]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[5]_net_1 ));
    OR2A \byte_ff_RNO[30]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_196)
        , .Y(\byte_ff_RNO[30]_net_1 ));
    MX2 \byte_ff_RNIOGIL[3]  (.A(\byte_ff[3]_net_1 ), .B(
        \buffer_ff[3]_net_1 ), .S(bypass_byte0), .Y(\crc_data_in0[3] ));
    OR2A \buffer_ff_RNO[17]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_287), .Y(\buffer_ff_RNO[17]_net_1 ));
    MX2 \crc_init_ff_RNO_0[7]  (.A(\crc_init_ff_3[7] ), .B(
        crc_init_out[7]), .S(un1_crc_init_en_1_0_net_1), .Y(N_138));
    DFN1 \byte_ff[28]  (.D(\byte_ff_RNO[28]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[28]_net_1 ));
    DFN1 \buffer_ff[15]  (.D(\buffer_ff_RNO[15]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[15]_net_1 ));
    MX2 \buffer_ff_RNO_0[7]  (.A(\buffer_ff[7]_net_1 ), .B(
        \bus_reversed[7] ), .S(buffer_en_0), .Y(N_277));
    NOR2B \crc_out_ff_RNO[10]  (.A(N_248), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[10]_net_1 ));
    MX2 \crc_init_ff_RNIMS9Q[23]  (.A(crc_init_out[23]), .B(
        \crc_out_ff[23]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[23] ));
    MX2 \crc_init_ff_RNIU28Q[18]  (.A(crc_init_out[18]), .B(
        \crc_out_ff[18]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[18] ));
    MX2 \crc_out_ff_RNO_0[20]  (.A(\crc_unit_out[20] ), .B(
        \crc_out_ff[20]_net_1 ), .S(state_byte_0[4]), .Y(N_258));
    OR2A \byte_ff_RNO[17]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_183)
        , .Y(\byte_ff_RNO[17]_net_1 ));
    MX2 \crc_init_ff_RNI05EL[9]  (.A(crc_init_out[9]), .B(
        \crc_out_ff[9]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[9] ));
    DFN1 \crc_poly_ff[11]  (.D(\crc_poly_ff_RNO[11]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[11]));
    NOR2 crc_poly_size_77_inst_1 (.A(crc_poly_size[1]), .B(
        crc_poly_size[0]), .Y(crc_poly_size_77));
    OR2A \byte_ff_RNO[22]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_188)
        , .Y(\byte_ff_RNO[22]_net_1 ));
    NOR2A crc_poly_size_75_0 (.A(crc_poly_size[1]), .B(
        crc_poly_size[0]), .Y(crc_poly_size_75_0_net_1));
    DFN1 \byte_ff[30]  (.D(\byte_ff_RNO[30]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[30]_net_1 ));
    DFN1 \buffer_ff[31]  (.D(\buffer_ff_RNO[31]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[31]_net_1 ));
    DFN1 \buffer_ff[14]  (.D(\buffer_ff_RNO[14]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[14]_net_1 ));
    DFN1 \crc_init_ff[24]  (.D(\crc_init_ff_RNO[24]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[24]));
    MX2 \crc_out_ff_RNO_0[3]  (.A(\crc_unit_out[3] ), .B(
        \crc_out_ff[3]_net_1 ), .S(state_byte[4]), .Y(N_241));
    MX2 \crc_init_ff_RNO_0[27]  (.A(\crc_init_ff_3[27] ), .B(
        crc_init_out[27]), .S(un1_crc_init_en_1_net_1), .Y(N_158));
    OR2A \crc_init_ff_RNO[10]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_141), .Y(\crc_init_ff_RNO[10]_net_1 ));
    OR2A \crc_init_ff_RNO_1[26]  (.A(crc_init_en), .B(N_332), .Y(
        \crc_init_ff_3[26] ));
    MX2 \buffer_ff_RNO_0[15]  (.A(\buffer_ff[15]_net_1 ), .B(
        \bus_reversed[15] ), .S(buffer_en_0), .Y(N_285));
    OR2A \buffer_ff_RNO[1]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_271), .Y(\buffer_ff_RNO[1]_net_1 ));
    MX2 \crc_out_ff_RNIB3HQ[13]  (.A(\crc_out_ff[18]_net_1 ), .B(
        \crc_out_ff[13]_net_1 ), .S(rev_out_type), .Y(crc_out[18]));
    DFN1 \crc_out_ff[27]  (.D(\crc_out_ff_RNO[27]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[27]_net_1 ));
    MX2 \crc_init_ff_RNO_0[11]  (.A(\crc_init_ff_3[11] ), .B(
        crc_init_out[11]), .S(un1_crc_init_en_1_0_net_1), .Y(N_142));
    MX2 \byte_ff_RNO_0[0]  (.A(\byte_ff[0]_net_1 ), .B(
        \buffer_ff[0]_net_1 ), .S(byte_en_0), .Y(N_166));
    OR2A \buffer_ff_RNO[7]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_277), .Y(\buffer_ff_RNO[7]_net_1 ));
    OR2A \crc_init_ff_RNO_1[16]  (.A(crc_init_en_0), .B(bus_wr_16), .Y(
        \crc_init_ff_3[16] ));
    MX2 \crc_init_ff_RNO_0[1]  (.A(\crc_init_ff_3[1] ), .B(
        crc_init_out[1]), .S(un1_crc_init_en_1_0_net_1), .Y(N_132));
    MX2 \crc_out_ff_RNI0QIL[11]  (.A(\crc_out_ff[11]_net_1 ), .B(
        \crc_out_ff[20]_net_1 ), .S(rev_out_type_0), .Y(crc_out[11]));
    MX2 \byte_ff_RNIQSRJ2[14]  (.A(N_110), .B(N_102), .S(N_294_0), .Y(
        \crc_data_in[6] ));
    DFN1 \crc_poly_ff[17]  (.D(\crc_poly_ff_RNO[17]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[17]));
    NOR2B \crc_idr_ff_RNO[0]  (.A(N_230), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_idr_ff_RNO[0]_net_1 ));
    MX2 \byte_ff_RNIV1SJ2[15]  (.A(N_111), .B(N_103), .S(N_294_0), .Y(
        \crc_data_in[7] ));
    MX2 \bf_size_ff_RNO_0[1]  (.A(\bf_size_ff[1]_net_1 ), .B(
        \bf_size_ff_4[1] ), .S(un1_buffer_en_net_1), .Y(N_164));
    OR2A \buffer_ff_RNO[21]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_291), .Y(\buffer_ff_RNO[21]_net_1 ));
    MX2 \crc_out_ff_RNIP47F[2]  (.A(\crc_out_ff[2]_net_1 ), .B(
        \crc_out_ff[29]_net_1 ), .S(rev_out_type_0), .Y(crc_out[2]));
    OR2A \crc_init_ff_RNO[0]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_131), .Y(\crc_init_ff_RNO[0]_net_1 ));
    DFN1 \crc_out_ff[8]  (.D(\crc_out_ff_RNO[8]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_out_ff[8]_net_1 ));
    DFN1 \crc_init_ff[8]  (.D(\crc_init_ff_RNO[8]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[8]));
    OR2A \crc_init_ff_RNO[5]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_136), .Y(\crc_init_ff_RNO[5]_net_1 ));
    MX2 \buffer_ff_RNO_0[0]  (.A(\buffer_ff[0]_net_1 ), .B(
        \bus_reversed[0] ), .S(buffer_en_0), .Y(N_270));
    OR2A \byte_ff_RNO[29]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_195)
        , .Y(\byte_ff_RNO[29]_net_1 ));
    NOR2B \crc_idr_ff_RNO[4]  (.A(N_234), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_idr_ff_RNO[4]_net_1 ));
    MX2 \crc_out_ff_RNO_0[1]  (.A(\crc_unit_out[1] ), .B(
        \crc_out_ff[1]_net_1 ), .S(state_byte[4]), .Y(N_239));
    OR2A \crc_init_ff_RNO_1[27]  (.A(crc_init_en), .B(N_333), .Y(
        \crc_init_ff_3[27] ));
    NOR2B \bf_size_ff_RNO[0]  (.A(N_163), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\bf_size_ff_RNO[0]_net_1 ));
    OR2A \crc_init_ff_RNO[13]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_144), .Y(\crc_init_ff_RNO[13]_net_1 ));
    DFN1 \byte_ff[22]  (.D(\byte_ff_RNO[22]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[22]_net_1 ));
    MX2 \crc_out_ff_RNIP47F[7]  (.A(\crc_out_ff[7]_net_1 ), .B(
        \crc_out_ff[24]_net_1 ), .S(rev_out_type_0), .Y(crc_out[7]));
    bit_reversal_32s_0_1_2_3_4s REV_IN (.rev_in_type_0({
        rev_in_type_0[0]}), .rev_in_type({rev_in_type[1], 
        rev_in_type[0]}), .bus_wr_0(bus_wr_0), .bus_wr_16(bus_wr_16), 
        .bus_wr_1(bus_wr_1), .bus_wr_25(bus_wr_25), .bus_wr_2(bus_wr_2)
        , .bus_wr_3(bus_wr_3), .bus_reversed({\bus_reversed[31] , 
        \bus_reversed[30] , \bus_reversed[29] , \bus_reversed[28] , 
        \bus_reversed[27] , \bus_reversed[26] , \bus_reversed[25] , 
        \bus_reversed[24] , \bus_reversed[23] , \bus_reversed[22] , 
        \bus_reversed[21] , \bus_reversed[20] , \bus_reversed[19] , 
        \bus_reversed[18] , \bus_reversed[17] , \bus_reversed[16] , 
        \bus_reversed[15] , \bus_reversed[14] , \bus_reversed[13] , 
        \bus_reversed[12] , \bus_reversed[11] , \bus_reversed[10] , 
        \bus_reversed[9] , \bus_reversed[8] , \bus_reversed[7] , 
        \bus_reversed[6] , \bus_reversed[5] , \bus_reversed[4] , 
        \bus_reversed[3] , \bus_reversed[2] , \bus_reversed[1] , 
        \bus_reversed[0] }), .N_358(N_358), .N_350(N_350), .N_351(
        N_351), .N_337(N_337), .N_366(N_366), .N_367(N_367), .N_357(
        N_357), .N_349(N_349), .N_352(N_352), .N_360(N_360), .N_336(
        N_336), .N_365(N_365), .N_356(N_356), .N_348(N_348), .N_353(
        N_353), .N_361(N_361), .N_335(N_335), .N_364(N_364), .N_332(
        N_332), .N_355(N_355), .N_362(N_362), .N_334(N_334), .N_333(
        N_333), .N_363(N_363), .N_347(N_347), .N_354(N_354));
    OR2A \crc_init_ff_RNO[16]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_147), .Y(\crc_init_ff_RNO[16]_net_1 ));
    OR2A \crc_poly_ff_RNO[8]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_206), .Y(\crc_poly_ff_RNO[8]_net_1 ));
    OR2A \byte_ff_RNO[15]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_181)
        , .Y(\byte_ff_RNO[15]_net_1 ));
    OR2A \crc_init_ff_RNO_1[17]  (.A(crc_init_en_0), .B(N_360), .Y(
        \crc_init_ff_3[17] ));
    MX2 \byte_ff_RNO_0[10]  (.A(\byte_ff[10]_net_1 ), .B(
        \buffer_ff[10]_net_1 ), .S(byte_en_0), .Y(N_176));
    MX2 \byte_ff_RNIMEIL[2]  (.A(\byte_ff[2]_net_1 ), .B(
        \buffer_ff[2]_net_1 ), .S(bypass_byte0), .Y(\crc_data_in0[2] ));
    MX2 \buffer_ff_RNO_0[3]  (.A(\buffer_ff[3]_net_1 ), .B(
        \bus_reversed[3] ), .S(buffer_en_0), .Y(N_273));
    NOR2B \crc_out_ff_RNO[24]  (.A(N_262), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[24]_net_1 ));
    DFN1 \crc_poly_ff[18]  (.D(\crc_poly_ff_RNO[18]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[18]));
    MX2 \crc_out_ff_RNIP47F[5]  (.A(\crc_out_ff[5]_net_1 ), .B(
        \crc_out_ff[26]_net_1 ), .S(rev_out_type_0), .Y(crc_out[5]));
    DFN1 \crc_poly_ff[24]  (.D(\crc_poly_ff_RNO[24]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[24]));
    OR2A \crc_init_ff_RNO_1[9]  (.A(crc_init_en), .B(N_352), .Y(
        \crc_init_ff_3[9] ));
    DFN1 \crc_poly_ff[13]  (.D(\crc_poly_ff_RNO[13]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[13]));
    MX2 \crc_idr_ff_RNO_0[3]  (.A(crc_idr_out[3]), .B(bus_wr_3), .S(
        crc_idr_en), .Y(N_233));
    MX2 \crc_init_ff_RNIMQDL[4]  (.A(crc_init_out[4]), .B(
        \crc_out_ff[4]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[4] ));
    OR2A \crc_poly_ff_RNO[1]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_199), .Y(\crc_poly_ff_RNO[1]_net_1 ));
    DFN1 \crc_init_ff[29]  (.D(\crc_init_ff_RNO[29]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[29]));
    NOR2B crc_poly_size_74_0 (.A(crc_poly_size[1]), .B(
        crc_poly_size[0]), .Y(crc_poly_size_74_0_net_1));
    MX2 \crc_poly_ff_RNO_0[25]  (.A(crc_poly_out[25]), .B(bus_wr_25), 
        .S(crc_poly_en_0), .Y(N_223));
    MX2 \crc_init_ff_RNIS08Q[17]  (.A(crc_init_out[17]), .B(
        \crc_out_ff[17]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[17] ));
    NOR2B \crc_out_ff_RNO[2]  (.A(N_240), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[2]_net_1 ));
    MX2 \crc_init_ff_RNIGK7Q[11]  (.A(crc_init_out[11]), .B(
        \crc_out_ff[11]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[11] ));
    DFN1 \crc_init_ff[26]  (.D(\crc_init_ff_RNO[26]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[26]));
    NOR2B \crc_poly_ff_RNO[6]  (.A(N_204), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[6]_net_1 ));
    OR2A \crc_init_ff_RNO_1[7]  (.A(crc_init_en), .B(N_350), .Y(
        \crc_init_ff_3[7] ));
    DFN1 \buffer_ff[25]  (.D(\buffer_ff_RNO[25]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[25]_net_1 ));
    DFN1 \crc_poly_ff[9]  (.D(\crc_poly_ff_RNO[9]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[9]));
    OR2A \crc_poly_ff_RNO[2]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_200), .Y(\crc_poly_ff_RNO[2]_net_1 ));
    MX2 \crc_idr_ff_RNO_0[0]  (.A(crc_idr_out[0]), .B(bus_wr_0), .S(
        crc_idr_en), .Y(N_230));
    OR2A un1_buffer_en (.A(N_56), .B(buffer_en), .Y(
        un1_buffer_en_net_1));
    OR2A \crc_init_ff_RNO[25]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_156), .Y(\crc_init_ff_RNO[25]_net_1 ));
    MX2 \crc_out_ff_RNIP47F[4]  (.A(\crc_out_ff[4]_net_1 ), .B(
        \crc_out_ff[27]_net_1 ), .S(rev_out_type_0), .Y(crc_out[4]));
    DFN1 \crc_idr_ff[2]  (.D(\crc_idr_ff_RNO[2]_net_1 ), .CLK(FAB_CLK), 
        .Q(crc_idr_out[2]));
    DFN1 \crc_init_ff[28]  (.D(\crc_init_ff_RNO[28]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[28]));
    OR2A \byte_ff_RNO[27]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_193)
        , .Y(\byte_ff_RNO[27]_net_1 ));
    OR2A \buffer_ff_RNO[31]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_301), .Y(\buffer_ff_RNO[31]_net_1 ));
    DFN1 \byte_ff[11]  (.D(\byte_ff_RNO[11]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[11]_net_1 ));
    MX2 \byte_ff_RNIUVQJ2[13]  (.A(N_109), .B(N_101), .S(N_294_0), .Y(
        \crc_data_in[5] ));
    NOR2B \crc_out_ff_RNO[9]  (.A(N_247), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[9]_net_1 ));
    DFN1 \buffer_ff[24]  (.D(\buffer_ff_RNO[24]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[24]_net_1 ));
    DFN1 \crc_init_ff[23]  (.D(\crc_init_ff_RNO[23]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[23]));
    MX2 \byte_ff_RNO_0[15]  (.A(\byte_ff[15]_net_1 ), .B(
        \buffer_ff[15]_net_1 ), .S(byte_en), .Y(N_181));
    MX2 \byte_ff_RNO_0[16]  (.A(\byte_ff[16]_net_1 ), .B(
        \buffer_ff[16]_net_1 ), .S(byte_en), .Y(N_182));
    MX2 \crc_out_ff_RNIP47F[8]  (.A(\crc_out_ff[8]_net_1 ), .B(
        \crc_out_ff[23]_net_1 ), .S(rev_out_type_0), .Y(crc_out[8]));
    OR2A \crc_init_ff_RNO_1[5]  (.A(crc_init_en), .B(N_348), .Y(
        \crc_init_ff_3[5] ));
    DFN1 \byte_ff[18]  (.D(\byte_ff_RNO[18]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[18]_net_1 ));
    OR2A \buffer_ff_RNO[18]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_288), .Y(\buffer_ff_RNO[18]_net_1 ));
    DFN1 \crc_init_ff[15]  (.D(\crc_init_ff_RNO[15]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[15]));
    DFN1 \crc_init_ff[5]  (.D(\crc_init_ff_RNO[5]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[5]));
    OR2A \byte_ff_RNO[1]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_167), 
        .Y(\byte_ff_RNO[1]_net_1 ));
    MX2 \crc_out_ff_RNIR56K[3]  (.A(\crc_out_ff[28]_net_1 ), .B(
        \crc_out_ff[3]_net_1 ), .S(rev_out_type), .Y(crc_out[28]));
    NOR2A un1_crc_init_en_1 (.A(N_56), .B(crc_init_en), .Y(
        un1_crc_init_en_1_net_1));
    OR2A \crc_init_ff_RNO[14]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_145), .Y(\crc_init_ff_RNO[14]_net_1 ));
    DFN1 \crc_poly_ff[26]  (.D(\crc_poly_ff_RNO[26]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[26]));
    MX2 \crc_init_ff_RNIIM7Q[12]  (.A(crc_init_out[12]), .B(
        \crc_out_ff[12]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[12] ));
    DFN1 \buffer_ff[10]  (.D(\buffer_ff_RNO[10]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[10]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[3]  (.A(crc_poly_out[3]), .B(bus_wr_3), .S(
        crc_poly_en), .Y(N_201));
    MX2 \byte_ff_RNICPAH2[9]  (.A(N_105), .B(N_97), .S(N_294_0), .Y(
        \crc_data_in[1] ));
    NOR2B \crc_out_ff_RNO[5]  (.A(N_243), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[5]_net_1 ));
    MX2 \crc_out_ff_RNIGS7F[0]  (.A(\crc_out_ff[0]_net_1 ), .B(
        \crc_out_ff[31]_net_1 ), .S(rev_out_type_0), .Y(crc_out[0]));
    MX2 \crc_init_ff_RNO_0[28]  (.A(\crc_init_ff_3[28] ), .B(
        crc_init_out[28]), .S(un1_crc_init_en_1_net_1), .Y(N_159));
    DFN1 \byte_ff[0]  (.D(\byte_ff_RNO[0]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[0]_net_1 ));
    MX2 \buffer_ff_RNO_0[2]  (.A(\buffer_ff[2]_net_1 ), .B(
        \bus_reversed[2] ), .S(buffer_en_0), .Y(N_272));
    OR2A \crc_init_ff_RNO[18]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_149), .Y(\crc_init_ff_RNO[18]_net_1 ));
    OR2A \buffer_ff_RNO[0]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_270), .Y(\buffer_ff_RNO[0]_net_1 ));
    OR2A \crc_poly_ff_RNO[10]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_208), .Y(\crc_poly_ff_RNO[10]_net_1 ));
    OR2A \buffer_ff_RNO[24]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_294), .Y(\buffer_ff_RNO[24]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[28]  (.A(crc_poly_out[28]), .B(N_334), .S(
        crc_poly_en), .Y(N_226));
    OR2A \byte_ff_RNO[25]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_191)
        , .Y(\byte_ff_RNO[25]_net_1 ));
    MX2 \buffer_ff_RNO_0[18]  (.A(\buffer_ff[18]_net_1 ), .B(
        \bus_reversed[18] ), .S(buffer_en), .Y(N_288));
    MX2 \crc_poly_ff_RNO_0[13]  (.A(crc_poly_out[13]), .B(N_356), .S(
        crc_poly_en_0), .Y(N_211));
    MX2 \crc_poly_ff_RNO_0[20]  (.A(crc_poly_out[20]), .B(N_363), .S(
        crc_poly_en_0), .Y(N_218));
    OR2A \crc_init_ff_RNO[12]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_143), .Y(\crc_init_ff_RNO[12]_net_1 ));
    MX2 \crc_init_ff_RNIMQ7Q[14]  (.A(crc_init_out[14]), .B(
        \crc_out_ff[14]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[14] ));
    MX2 \byte_ff_RNO_0[24]  (.A(\byte_ff[24]_net_1 ), .B(
        \buffer_ff[24]_net_1 ), .S(byte_en), .Y(N_190));
    MX2 \crc_idr_ff_RNO_0[6]  (.A(crc_idr_out[6]), .B(N_349), .S(
        crc_idr_en), .Y(N_236));
    OR2A \crc_init_ff_RNO[1]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_132), .Y(\crc_init_ff_RNO[1]_net_1 ));
    OR2A \crc_init_ff_RNO_1[28]  (.A(crc_init_en), .B(N_334), .Y(
        \crc_init_ff_3[28] ));
    DFN1 \byte_ff[12]  (.D(\byte_ff_RNO[12]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[12]_net_1 ));
    OR2A \buffer_ff_RNO[8]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_278), .Y(\buffer_ff_RNO[8]_net_1 ));
    NOR2B \crc_out_ff_RNO[23]  (.A(N_261), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[23]_net_1 ));
    OR2A \crc_init_ff_RNO_1[0]  (.A(crc_init_en), .B(bus_wr_0), .Y(
        \crc_init_ff_3[0] ));
    DFN1 \crc_out_ff[9]  (.D(\crc_out_ff_RNO[9]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_out_ff[9]_net_1 ));
    MX2 \crc_init_ff_RNIIMDL[2]  (.A(crc_init_out[2]), .B(
        \crc_out_ff[2]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[2] ));
    OR2A \crc_init_ff_RNO_1[18]  (.A(crc_init_en_0), .B(N_361), .Y(
        \crc_init_ff_3[18] ));
    DFN1 \crc_idr_ff[3]  (.D(\crc_idr_ff_RNO[3]_net_1 ), .CLK(FAB_CLK), 
        .Q(crc_idr_out[3]));
    MX2 \crc_poly_ff_RNO_0[29]  (.A(crc_poly_out[29]), .B(N_335), .S(
        crc_poly_en), .Y(N_227));
    DFN1 \crc_out_ff[14]  (.D(\crc_out_ff_RNO[14]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[14]_net_1 ));
    NOR2B \crc_poly_ff_RNO[17]  (.A(N_215), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[17]_net_1 ));
    MX2 \crc_idr_ff_RNO_0[7]  (.A(crc_idr_out[7]), .B(N_350), .S(
        crc_idr_en), .Y(N_237));
    NOR2B crc_init_sel_ff_RNI2BI2B (.A(N_165), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(
        crc_init_sel_ff_RNI2BI2B_net_1));
    MX2 \byte_ff_RNI07BA1[23]  (.A(\byte_ff[23]_net_1 ), .B(
        \crc_data_in0[7] ), .S(N_128), .Y(N_103));
    NOR2B \crc_out_ff_RNO[16]  (.A(N_254), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[16]_net_1 ));
    MX2 \crc_out_ff_RNO_0[26]  (.A(\crc_unit_out[26] ), .B(
        \crc_out_ff[26]_net_1 ), .S(state_byte[4]), .Y(N_264));
    MX2 \byte_ff_RNO_0[2]  (.A(\byte_ff[2]_net_1 ), .B(
        \buffer_ff[2]_net_1 ), .S(byte_en_0), .Y(N_168));
    DFN1 \crc_poly_ff[6]  (.D(\crc_poly_ff_RNO[6]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[6]));
    NOR2B \crc_out_ff_RNO[1]  (.A(N_239), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[1]_net_1 ));
    NOR2B \crc_poly_ff_RNO[20]  (.A(N_218), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[20]_net_1 ));
    DFN1 \crc_idr_ff[5]  (.D(\crc_idr_ff_RNO[5]_net_1 ), .CLK(FAB_CLK), 
        .Q(crc_idr_out[5]));
    NOR2B \crc_out_ff_RNO[20]  (.A(N_258), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[20]_net_1 ));
    MX2 \crc_out_ff_RNIP47F[9]  (.A(\crc_out_ff[9]_net_1 ), .B(
        \crc_out_ff[22]_net_1 ), .S(rev_out_type_0), .Y(crc_out[9]));
    MX2 \crc_out_ff_RNO_0[25]  (.A(\crc_unit_out[25] ), .B(
        \crc_out_ff[25]_net_1 ), .S(state_byte_0[4]), .Y(N_263));
    MX2 \crc_out_ff_RNI92IL_0[15]  (.A(\crc_out_ff[15]_net_1 ), .B(
        \crc_out_ff[16]_net_1 ), .S(rev_out_type_0), .Y(crc_out[15]));
    DFN1 \crc_out_ff[1]  (.D(\crc_out_ff_RNO[1]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_out_ff[1]_net_1 ));
    DFN1 \byte_ff[3]  (.D(\byte_ff_RNO[3]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[3]_net_1 ));
    MX2 \crc_init_ff_RNIIO9Q[21]  (.A(crc_init_out[21]), .B(
        \crc_out_ff[21]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[21] ));
    MX2 \byte_ff_RNISKIL[5]  (.A(\byte_ff[5]_net_1 ), .B(
        \buffer_ff[5]_net_1 ), .S(bypass_byte0), .Y(\crc_data_in0[5] ));
    MX2 \size_ff_RNI7H3P[1]  (.A(\size_ff[1]_net_1 ), .B(
        \bf_size_ff[1]_net_1 ), .S(N_118_1), .Y(size_in[1]));
    OR2A \byte_ff_RNO[9]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_175), 
        .Y(\byte_ff_RNO[9]_net_1 ));
    DFN1 \byte_ff[8]  (.D(\byte_ff_RNO[8]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[8]_net_1 ));
    OR2A \crc_init_ff_RNO_1[8]  (.A(crc_init_en), .B(N_351), .Y(
        \crc_init_ff_3[8] ));
    MX2 \crc_init_ff_RNO_0[16]  (.A(\crc_init_ff_3[16] ), .B(
        crc_init_out[16]), .S(un1_crc_init_en_1_net_1), .Y(N_147));
    MX2 \crc_out_ff_RNO_0[14]  (.A(\crc_unit_out[14] ), .B(
        \crc_out_ff[14]_net_1 ), .S(state_byte_0[4]), .Y(N_252));
    DFN1 \buffer_ff[20]  (.D(\buffer_ff_RNO[20]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[20]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[26]  (.A(crc_poly_out[26]), .B(N_332), .S(
        crc_poly_en), .Y(N_224));
    MX2 \crc_out_ff_RNIR56K[2]  (.A(\crc_out_ff[29]_net_1 ), .B(
        \crc_out_ff[2]_net_1 ), .S(rev_out_type), .Y(crc_out[29]));
    MX2 \crc_idr_ff_RNO_0[2]  (.A(crc_idr_out[2]), .B(bus_wr_2), .S(
        crc_idr_en), .Y(N_232));
    OR2A \crc_poly_ff_RNO[7]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_205), .Y(\crc_poly_ff_RNO[7]_net_1 ));
    MX2 \crc_init_ff_RNI00UR[27]  (.A(crc_init_out[27]), .B(
        \crc_out_ff[27]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[27] ));
    DFN1 \crc_poly_ff[14]  (.D(\crc_poly_ff_RNO[14]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[14]));
    MX2 \crc_init_ff_RNO_0[23]  (.A(\crc_init_ff_3[23] ), .B(
        crc_init_out[23]), .S(un1_crc_init_en_1_net_1), .Y(N_154));
    MX2 \byte_ff_RNO_0[6]  (.A(\byte_ff[6]_net_1 ), .B(
        \buffer_ff[6]_net_1 ), .S(byte_en_0), .Y(N_172));
    DFN1 \buffer_ff[8]  (.D(\buffer_ff_RNO[8]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[8]_net_1 ));
    NOR2B \crc_poly_ff_RNO[27]  (.A(N_225), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[27]_net_1 ));
    DFN1 \buffer_ff[18]  (.D(\buffer_ff_RNO[18]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[18]_net_1 ));
    OR2A \crc_init_ff_RNO[27]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_158), .Y(\crc_init_ff_RNO[27]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[11]  (.A(crc_poly_out[11]), .B(N_354), .S(
        crc_poly_en_0), .Y(N_209));
    DFN1 \crc_init_ff[0]  (.D(\crc_init_ff_RNO[0]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[0]));
    NOR2B \crc_poly_ff_RNO[15]  (.A(N_213), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[15]_net_1 ));
    MX2 \byte_ff_RNIQV9A1[18]  (.A(\byte_ff[18]_net_1 ), .B(
        \crc_data_in0[2] ), .S(N_128), .Y(N_98));
    DFN1 \crc_init_ff[10]  (.D(\crc_init_ff_RNO[10]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[10]));
    MX2 \byte_ff_RNINTAA1[20]  (.A(\byte_ff[20]_net_1 ), .B(
        \crc_data_in0[4] ), .S(N_128), .Y(N_100));
    DFN1 \buffer_ff[4]  (.D(\buffer_ff_RNO[4]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[4]_net_1 ));
    OR2A \crc_init_ff_RNO[3]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_134), .Y(\crc_init_ff_RNO[3]_net_1 ));
    MX2 \crc_init_ff_RNO_0[25]  (.A(\crc_init_ff_3[25] ), .B(
        crc_init_out[25]), .S(un1_crc_init_en_1_net_1), .Y(N_156));
    MX2 \byte_ff_RNI69AP[12]  (.A(\byte_ff[28]_net_1 ), .B(
        \byte_ff[12]_net_1 ), .S(N_128), .Y(N_108));
    DFN1 \crc_poly_ff[2]  (.D(\crc_poly_ff_RNO[2]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[2]));
    MX2 \buffer_ff_RNO_0[25]  (.A(\buffer_ff[25]_net_1 ), .B(
        \bus_reversed[25] ), .S(buffer_en), .Y(N_295));
    MX2 \byte_ff_RNIT2AA1[19]  (.A(\byte_ff[19]_net_1 ), .B(
        \crc_data_in0[3] ), .S(N_128), .Y(N_99));
    MX2 \crc_init_ff_RNO_0[17]  (.A(\crc_init_ff_3[17] ), .B(
        crc_init_out[17]), .S(un1_crc_init_en_1_net_1), .Y(N_148));
    MX2 \crc_poly_ff_RNO_0[22]  (.A(crc_poly_out[22]), .B(N_365), .S(
        crc_poly_en_0), .Y(N_220));
    NOR2B \crc_out_ff_RNO[11]  (.A(N_249), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[11]_net_1 ));
    DFN1 \crc_init_ff[30]  (.D(\crc_init_ff_RNO[30]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[30]));
    OR2A \buffer_ff_RNO[11]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_281), .Y(\buffer_ff_RNO[11]_net_1 ));
    DFN1 \crc_poly_ff[30]  (.D(\crc_poly_ff_RNO[30]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[30]));
    DFN1 \crc_init_ff[1]  (.D(\crc_init_ff_RNO[1]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[1]));
    DFN1 \byte_ff[31]  (.D(\byte_ff_RNO[31]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[31]_net_1 ));
    MX2 \crc_out_ff_RNI2RHQ[10]  (.A(\crc_out_ff[21]_net_1 ), .B(
        \crc_out_ff[10]_net_1 ), .S(rev_out_type), .Y(crc_out[21]));
    MX2 \crc_out_ff_RNI92IL[15]  (.A(\crc_out_ff[16]_net_1 ), .B(
        \crc_out_ff[15]_net_1 ), .S(rev_out_type_0), .Y(crc_out[16]));
    OR2A \crc_init_ff_RNO_1[6]  (.A(crc_init_en), .B(N_349), .Y(
        \crc_init_ff_3[6] ));
    DFN1 \buffer_ff[16]  (.D(\buffer_ff_RNO[16]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[16]_net_1 ));
    DFN1 \crc_init_ff[7]  (.D(\crc_init_ff_RNO[7]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[7]));
    MX2 \buffer_ff_RNO_0[17]  (.A(\buffer_ff[17]_net_1 ), .B(
        \bus_reversed[17] ), .S(buffer_en_0), .Y(N_287));
    MX2 \byte_ff_RNIQ0BA1[21]  (.A(\byte_ff[21]_net_1 ), .B(
        \crc_data_in0[5] ), .S(N_128), .Y(N_101));
    MX2 \crc_init_ff_RNI058Q[19]  (.A(crc_init_out[19]), .B(
        \crc_out_ff[19]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[19] ));
    MX2 \crc_out_ff_RNIP47F[6]  (.A(\crc_out_ff[6]_net_1 ), .B(
        \crc_out_ff[25]_net_1 ), .S(rev_out_type_0), .Y(crc_out[6]));
    OR2A \crc_init_ff_RNO_1[23]  (.A(crc_init_en_0), .B(N_366), .Y(
        \crc_init_ff_3[23] ));
    MX2 \crc_init_ff_RNO_0[6]  (.A(\crc_init_ff_3[6] ), .B(
        crc_init_out[6]), .S(un1_crc_init_en_1_0_net_1), .Y(N_137));
    OR2A \byte_ff_RNO[5]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_171), 
        .Y(\byte_ff_RNO[5]_net_1 ));
    MX2 \crc_out_ff_RNO_0[13]  (.A(\crc_unit_out[13] ), .B(
        \crc_out_ff[13]_net_1 ), .S(state_byte_0[4]), .Y(N_251));
    OR2A \buffer_ff_RNO[4]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_274), .Y(\buffer_ff_RNO[4]_net_1 ));
    DFN1 \byte_ff[1]  (.D(\byte_ff_RNO[1]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[1]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[0]  (.A(crc_poly_out[0]), .B(bus_wr_0), .S(
        crc_poly_en), .Y(N_198));
    OR2A \crc_init_ff_RNO[6]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_137), .Y(\crc_init_ff_RNO[6]_net_1 ));
    OR2A \crc_init_ff_RNO_1[13]  (.A(crc_init_en_0), .B(N_356), .Y(
        \crc_init_ff_3[13] ));
    MX2 \buffer_ff_RNO_0[6]  (.A(\buffer_ff[6]_net_1 ), .B(
        \bus_reversed[6] ), .S(buffer_en_0), .Y(N_276));
    OR2A \crc_init_ff_RNO_1[25]  (.A(crc_init_en_0), .B(bus_wr_25), .Y(
        \crc_init_ff_3[25] ));
    NOR2A un1_crc_init_en_1_0 (.A(N_56), .B(crc_init_en), .Y(
        un1_crc_init_en_1_0_net_1));
    MX2 \crc_poly_ff_RNO_0[24]  (.A(crc_poly_out[24]), .B(N_367), .S(
        crc_poly_en_0), .Y(N_222));
    MX2 \size_ff_RNO_0[0]  (.A(\size_ff[0]_net_1 ), .B(
        \bf_size_ff[0]_net_1 ), .S(byte_en_0), .Y(N_129));
    MX2 \crc_poly_ff_RNO_0[5]  (.A(crc_poly_out[5]), .B(N_348), .S(
        crc_poly_en), .Y(N_203));
    MX2 \crc_out_ff_RNO_0[4]  (.A(\crc_unit_out[4] ), .B(
        \crc_out_ff[4]_net_1 ), .S(state_byte[4]), .Y(N_242));
    OR2A \buffer_ff_RNO[26]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_296), .Y(\buffer_ff_RNO[26]_net_1 ));
    NOR2B \crc_poly_ff_RNO[18]  (.A(N_216), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[18]_net_1 ));
    MX2 \buffer_ff_RNO_0[13]  (.A(\buffer_ff[13]_net_1 ), .B(
        \bus_reversed[13] ), .S(buffer_en_0), .Y(N_283));
    OR2A \crc_init_ff_RNO_1[15]  (.A(crc_init_en_0), .B(N_358), .Y(
        \crc_init_ff_3[15] ));
    MX2 \crc_out_ff_RNO_0[2]  (.A(\crc_unit_out[2] ), .B(
        \crc_out_ff[2]_net_1 ), .S(state_byte[4]), .Y(N_240));
    MX2 \crc_out_ff_RNIB3HQ[14]  (.A(\crc_out_ff[17]_net_1 ), .B(
        \crc_out_ff[14]_net_1 ), .S(rev_out_type), .Y(crc_out[17]));
    MX2 \byte_ff_RNO_0[14]  (.A(\byte_ff[14]_net_1 ), .B(
        \buffer_ff[14]_net_1 ), .S(byte_en_0), .Y(N_180));
    DFN1 \buffer_ff[13]  (.D(\buffer_ff_RNO[13]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[13]_net_1 ));
    OR2A \buffer_ff_RNO[25]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_295), .Y(\buffer_ff_RNO[25]_net_1 ));
    NOR2B \crc_out_ff_RNO[0]  (.A(N_238), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[0]_net_1 ));
    OR2A \buffer_ff_RNO[23]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_293), .Y(\buffer_ff_RNO[23]_net_1 ));
    NOR2B \crc_poly_ff_RNO[25]  (.A(N_223), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[25]_net_1 ));
    MX2 \crc_out_ff_RNI92IL[14]  (.A(\crc_out_ff[14]_net_1 ), .B(
        \crc_out_ff[17]_net_1 ), .S(rev_out_type_0), .Y(crc_out[14]));
    DFN1 \crc_poly_ff[16]  (.D(\crc_poly_ff_RNO[16]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[16]));
    OR2A \byte_ff_RNO[7]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_173), 
        .Y(\byte_ff_RNO[7]_net_1 ));
    DFN1 crc_init_sel_ff_0_0 (.D(crc_init_sel_ff_RNI2BI2B_net_1), .CLK(
        FAB_CLK), .Q(crc_init_sel_ff_0));
    MX2 \crc_out_ff_RNI92IL[13]  (.A(\crc_out_ff[13]_net_1 ), .B(
        \crc_out_ff[18]_net_1 ), .S(rev_out_type_0), .Y(crc_out[13]));
    OR2A \buffer_ff_RNO[22]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_292), .Y(\buffer_ff_RNO[22]_net_1 ));
    DFN1 \crc_out_ff[30]  (.D(\crc_out_ff_RNO[30]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[30]_net_1 ));
    DFN1 \crc_init_ff[4]  (.D(\crc_init_ff_RNO[4]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[4]));
    DFN1 \crc_out_ff[31]  (.D(\crc_out_ff_RNO[31]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[31]_net_1 ));
    MX2 \crc_out_ff_RNO_0[21]  (.A(\crc_unit_out[21] ), .B(
        \crc_out_ff[21]_net_1 ), .S(state_byte_0[4]), .Y(N_259));
    DFN1 \crc_poly_ff[4]  (.D(\crc_poly_ff_RNO[4]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[4]));
    NOR2B \crc_idr_ff_RNO[1]  (.A(N_231), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_idr_ff_RNO[1]_net_1 ));
    MX2 \crc_init_ff_RNIGM9Q[20]  (.A(crc_init_out[20]), .B(
        \crc_out_ff[20]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[20] ));
    DFN1 \crc_init_ff[12]  (.D(\crc_init_ff_RNO[12]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[12]));
    OR2A \byte_ff_RNO[8]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_174), 
        .Y(\byte_ff_RNO[8]_net_1 ));
    OR2A \crc_init_ff_RNO[4]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_135), .Y(\crc_init_ff_RNO[4]_net_1 ));
    OR2A \crc_init_ff_RNO[7]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_138), .Y(\crc_init_ff_RNO[7]_net_1 ));
    MX2 \crc_out_ff_RNIR56K[5]  (.A(\crc_out_ff[26]_net_1 ), .B(
        \crc_out_ff[5]_net_1 ), .S(rev_out_type), .Y(crc_out[26]));
    MX2 \crc_init_ff_RNO_0[3]  (.A(\crc_init_ff_3[3] ), .B(
        crc_init_out[3]), .S(un1_crc_init_en_1_0_net_1), .Y(N_134));
    NOR2B \size_ff_RNO[0]  (.A(N_129), .B(crc_ahb_ip_MSS_0_M2F_RESET_N)
        , .Y(\size_ff_RNO[0]_net_1 ));
    DFN1 \buffer_ff[30]  (.D(\buffer_ff_RNO[30]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[30]_net_1 ));
    DFN1 \crc_idr_ff[4]  (.D(\crc_idr_ff_RNO[4]_net_1 ), .CLK(FAB_CLK), 
        .Q(crc_idr_out[4]));
    DFN1 \crc_poly_ff[8]  (.D(\crc_poly_ff_RNO[8]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[8]));
    DFN1 \crc_poly_ff[22]  (.D(\crc_poly_ff_RNO[22]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[22]));
    OR2A \bf_size_ff_RNO_1[1]  (.A(buffer_en), .B(bus_size[1]), .Y(
        \bf_size_ff_4[1] ));
    DFN1 \crc_init_ff[11]  (.D(\crc_init_ff_RNO[11]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[11]));
    NOR2B \crc_idr_ff_RNO[6]  (.A(N_236), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_idr_ff_RNO[6]_net_1 ));
    MX2 \byte_ff_RNI37BP[15]  (.A(\byte_ff[31]_net_1 ), .B(
        \byte_ff[15]_net_1 ), .S(N_128), .Y(N_111));
    MX2 \byte_ff_RNI25AP[10]  (.A(\byte_ff[26]_net_1 ), .B(
        \byte_ff[10]_net_1 ), .S(N_128), .Y(N_106));
    DFN1 \buffer_ff[28]  (.D(\buffer_ff_RNO[28]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[28]_net_1 ));
    DFN1 \crc_init_ff[31]  (.D(\crc_init_ff_RNO[31]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[31]));
    NOR2B \crc_poly_ff_RNO[3]  (.A(N_201), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[3]_net_1 ));
    DFN1 \byte_ff[9]  (.D(\byte_ff_RNO[9]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[9]_net_1 ));
    NOR2B \crc_poly_ff_RNO[28]  (.A(N_226), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[28]_net_1 ));
    MX2 \crc_init_ff_RNIEI7Q[10]  (.A(crc_init_out[10]), .B(
        \crc_out_ff[10]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[10] ));
    DFN1 \buffer_ff[3]  (.D(\buffer_ff_RNO[3]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[3]_net_1 ));
    MX2 \crc_init_ff_RNO_0[5]  (.A(\crc_init_ff_3[5] ), .B(
        crc_init_out[5]), .S(un1_crc_init_en_1_0_net_1), .Y(N_136));
    DFN1 \crc_init_ff[17]  (.D(\crc_init_ff_RNO[17]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[17]));
    OR2A \byte_ff_RNO[31]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_197)
        , .Y(\byte_ff_RNO[31]_net_1 ));
    MX2 \crc_init_ff_RNO_0[4]  (.A(\crc_init_ff_3[4] ), .B(
        crc_init_out[4]), .S(un1_crc_init_en_1_0_net_1), .Y(N_135));
    DFN1 \buffer_ff[26]  (.D(\buffer_ff_RNO[26]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[26]_net_1 ));
    NOR2A crc_poly_size_76 (.A(crc_poly_size[0]), .B(crc_poly_size[1]), 
        .Y(crc_poly_size_76_net_1));
    NOR2B \crc_out_ff_RNO[18]  (.A(N_256), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[18]_net_1 ));
    MX2 \crc_out_ff_RNO_0[29]  (.A(\crc_unit_out[29] ), .B(
        \crc_out_ff[29]_net_1 ), .S(state_byte[4]), .Y(N_267));
    MX2 \crc_out_ff_RNO_0[28]  (.A(\crc_unit_out[28] ), .B(
        \crc_out_ff[28]_net_1 ), .S(state_byte[4]), .Y(N_266));
    MX2 \crc_out_ff_RNO_0[17]  (.A(\crc_unit_out[17] ), .B(
        \crc_out_ff[17]_net_1 ), .S(state_byte_0[4]), .Y(N_255));
    MX2 \byte_ff_RNO_0[3]  (.A(\byte_ff[3]_net_1 ), .B(
        \buffer_ff[3]_net_1 ), .S(byte_en_0), .Y(N_169));
    OR2A \byte_ff_RNO[10]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_176)
        , .Y(\byte_ff_RNO[10]_net_1 ));
    MX2 \byte_ff_RNI8BAP[13]  (.A(\byte_ff[29]_net_1 ), .B(
        \byte_ff[13]_net_1 ), .S(N_128), .Y(N_109));
    OR2A \crc_init_ff_RNO[29]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_160), .Y(\crc_init_ff_RNO[29]_net_1 ));
    OR2A \buffer_ff_RNO[14]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_284), .Y(\buffer_ff_RNO[14]_net_1 ));
    MX2 \crc_poly_ff_RNO_0[31]  (.A(crc_poly_out[31]), .B(N_337), .S(
        crc_poly_en), .Y(N_229));
    MX2 \buffer_ff_RNO_0[10]  (.A(\buffer_ff[10]_net_1 ), .B(
        \bus_reversed[10] ), .S(buffer_en_0), .Y(N_280));
    OR2A \crc_poly_ff_RNO[4]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_202), .Y(\crc_poly_ff_RNO[4]_net_1 ));
    MX2 \byte_ff_RNO_0[21]  (.A(\byte_ff[21]_net_1 ), .B(
        \buffer_ff[21]_net_1 ), .S(byte_en), .Y(N_187));
    DFN1 \crc_out_ff[10]  (.D(\crc_out_ff_RNO[10]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[10]_net_1 ));
    DFN1 \crc_out_ff[11]  (.D(\crc_out_ff_RNO[11]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[11]_net_1 ));
    MX2 \crc_out_ff_RNO_0[12]  (.A(\crc_unit_out[12] ), .B(
        \crc_out_ff[12]_net_1 ), .S(state_byte_0[4]), .Y(N_250));
    MX2 \crc_init_ff_RNO_0[18]  (.A(\crc_init_ff_3[18] ), .B(
        crc_init_out[18]), .S(un1_crc_init_en_1_net_1), .Y(N_149));
    MX2 \crc_init_ff_RNIMNVR[31]  (.A(crc_init_out[31]), .B(
        \crc_out_ff[31]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[31] ));
    DFN1 \buffer_ff[1]  (.D(\buffer_ff_RNO[1]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[1]_net_1 ));
    MX2 \byte_ff_RNO_0[30]  (.A(\byte_ff[30]_net_1 ), .B(
        \buffer_ff[30]_net_1 ), .S(byte_en), .Y(N_196));
    crc_parallel_32s_8s_4294967295_0 CRC_UNIT (.crc_poly_out({
        crc_poly_out[31], crc_poly_out[30], crc_poly_out[29], 
        crc_poly_out[28], crc_poly_out[27], crc_poly_out[26], 
        crc_poly_out[25], crc_poly_out[24], crc_poly_out[23], 
        crc_poly_out[22], crc_poly_out[21], crc_poly_out[20], 
        crc_poly_out[19], crc_poly_out[18], crc_poly_out[17], 
        crc_poly_out[16], crc_poly_out[15], crc_poly_out[14], 
        crc_poly_out[13], crc_poly_out[12], crc_poly_out[11], 
        crc_poly_out[10], crc_poly_out[9], crc_poly_out[8], 
        crc_poly_out[7], crc_poly_out[6], crc_poly_out[5], 
        crc_poly_out[4], crc_poly_out[3], crc_poly_out[2], 
        crc_poly_out[1], crc_poly_out[0]}), .crc_init_mux({
        \crc_init_mux[31] , \crc_init_mux[30] , \crc_init_mux[29] , 
        \crc_init_mux[28] , \crc_init_mux[27] , \crc_init_mux[26] , 
        \crc_init_mux[25] , \crc_init_mux[24] , \crc_init_mux[23] , 
        \crc_init_mux[22] , \crc_init_mux[21] , \crc_init_mux[20] , 
        \crc_init_mux[19] , \crc_init_mux[18] , \crc_init_mux[17] , 
        \crc_init_mux[16] , \crc_init_mux[15] , \crc_init_mux[14] , 
        \crc_init_mux[13] , \crc_init_mux[12] , \crc_init_mux[11] , 
        \crc_init_mux[10] , \crc_init_mux[9] , \crc_init_mux[8] , 
        \crc_init_mux[7] , \crc_init_mux[6] , \crc_init_mux[5] , 
        \crc_init_mux[4] , \crc_init_mux[3] , \crc_init_mux[2] , 
        \crc_init_mux[1] , \crc_init_mux[0] }), .crc_data_in({
        \crc_data_in[7] , \crc_data_in[6] , \crc_data_in[5] , 
        \crc_data_in[4] , \crc_data_in[3] , \crc_data_in[2] , 
        \crc_data_in[1] , \crc_data_in[0] }), .crc_unit_out({
        \crc_unit_out[31] , \crc_unit_out[30] , \crc_unit_out[29] , 
        \crc_unit_out[28] , \crc_unit_out[27] , \crc_unit_out[26] , 
        \crc_unit_out[25] , \crc_unit_out[24] , \crc_unit_out[23] , 
        \crc_unit_out[22] , \crc_unit_out[21] , \crc_unit_out[20] , 
        \crc_unit_out[19] , \crc_unit_out[18] , \crc_unit_out[17] , 
        \crc_unit_out[16] , \crc_unit_out[15] , \crc_unit_out[14] , 
        \crc_unit_out[13] , \crc_unit_out[12] , \crc_unit_out[11] , 
        \crc_unit_out[10] , \crc_unit_out[9] , \crc_unit_out[8] , 
        \crc_unit_out[7] , \crc_unit_out[6] , \crc_unit_out[5] , 
        \crc_unit_out[4] , \crc_unit_out[3] , \crc_unit_out[2] , 
        \crc_unit_out[1] , \crc_unit_out[0] }), .crc_poly_size_76(
        crc_poly_size_76_net_1), .crc_poly_size_77(crc_poly_size_77_0), 
        .crc_poly_size_74(crc_poly_size_74_net_1), .crc_poly_size_75_0(
        crc_poly_size_75_0_net_1), .crc_poly_size_76_0(
        crc_poly_size_76_0_net_1), .crc_poly_size_74_0(
        crc_poly_size_74_0_net_1), .crc_poly_size_76_1(
        crc_poly_size_76_1_net_1), .crc_poly_size_75(
        crc_poly_size_75_net_1));
    MX2 \crc_out_ff_RNO_0[30]  (.A(\crc_unit_out[30] ), .B(
        \crc_out_ff[30]_net_1 ), .S(state_byte[4]), .Y(N_268));
    MX2 \buffer_ff_RNO_0[28]  (.A(\buffer_ff[28]_net_1 ), .B(
        \bus_reversed[28] ), .S(buffer_en), .Y(N_298));
    DFN1 \buffer_ff[23]  (.D(\buffer_ff_RNO[23]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[23]_net_1 ));
    MX2 \crc_idr_ff_RNO_0[5]  (.A(crc_idr_out[5]), .B(N_348), .S(
        crc_idr_en), .Y(N_235));
    DFN1 \crc_out_ff[12]  (.D(\crc_out_ff_RNO[12]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[12]_net_1 ));
    DFN1 \crc_init_ff[2]  (.D(\crc_init_ff_RNO[2]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[2]));
    DFN1 \crc_idr_ff[1]  (.D(\crc_idr_ff_RNO[1]_net_1 ), .CLK(FAB_CLK), 
        .Q(crc_idr_out[1]));
    MX2 \byte_ff_RNO_0[28]  (.A(\byte_ff[28]_net_1 ), .B(
        \buffer_ff[28]_net_1 ), .S(byte_en), .Y(N_194));
    OR2A \buffer_ff_RNO[6]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_276), .Y(\buffer_ff_RNO[6]_net_1 ));
    NOR2B \crc_out_ff_RNO[26]  (.A(N_264), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[26]_net_1 ));
    DFN1 \crc_init_ff[14]  (.D(\crc_init_ff_RNO[14]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[14]));
    VCC VCC_i (.Y(VCC));
    DFN1 \crc_out_ff[16]  (.D(\crc_out_ff_RNO[16]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[16]_net_1 ));
    DFN1 \crc_idr_ff[7]  (.D(\crc_idr_ff_RNO[7]_net_1 ), .CLK(FAB_CLK), 
        .Q(crc_idr_out[7]));
    MX2 \crc_init_ff_RNIOS7Q[15]  (.A(crc_init_out[15]), .B(
        \crc_out_ff[15]_net_1 ), .S(crc_init_sel_ff_0), .Y(
        \crc_init_mux[15] ));
    MX2 \crc_poly_ff_RNO_0[9]  (.A(crc_poly_out[9]), .B(N_352), .S(
        crc_poly_en), .Y(N_207));
    MX2 \byte_ff_RNIPQQJ2[12]  (.A(N_108), .B(N_100), .S(N_294_0), .Y(
        \crc_data_in[4] ));
    DFN1 \size_ff[0]  (.D(\size_ff_RNO[0]_net_1 ), .CLK(FAB_CLK), .Q(
        \size_ff[0]_net_1 ));
    OR2A \byte_ff_RNO[14]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(N_180)
        , .Y(\byte_ff_RNO[14]_net_1 ));
    DFN1 \crc_out_ff[24]  (.D(\crc_out_ff_RNO[24]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[24]_net_1 ));
    NOR2A crc_poly_size_76_0 (.A(crc_poly_size[0]), .B(
        crc_poly_size[1]), .Y(crc_poly_size_76_0_net_1));
    MX2 \crc_init_ff_RNO_0[20]  (.A(\crc_init_ff_3[20] ), .B(
        crc_init_out[20]), .S(un1_crc_init_en_1_net_1), .Y(N_151));
    DFN1 \byte_ff[26]  (.D(\byte_ff_RNO[26]_net_1 ), .CLK(FAB_CLK), .Q(
        \byte_ff[26]_net_1 ));
    MX2 \crc_out_ff_RNIR56K[4]  (.A(\crc_out_ff[27]_net_1 ), .B(
        \crc_out_ff[4]_net_1 ), .S(rev_out_type), .Y(crc_out[27]));
    NOR2B \crc_out_ff_RNO[15]  (.A(N_253), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[15]_net_1 ));
    MX2 \crc_init_ff_RNIQUDL[6]  (.A(crc_init_out[6]), .B(
        \crc_out_ff[6]_net_1 ), .S(crc_init_sel_ff_net_1), .Y(
        \crc_init_mux[6] ));
    NOR2B \crc_out_ff_RNO[30]  (.A(N_268), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[30]_net_1 ));
    DFN1 \crc_out_ff[18]  (.D(\crc_out_ff_RNO[18]_net_1 ), .CLK(
        FAB_CLK), .Q(\crc_out_ff[18]_net_1 ));
    MX2 \buffer_ff_RNO_0[11]  (.A(\buffer_ff[11]_net_1 ), .B(
        \bus_reversed[11] ), .S(buffer_en_0), .Y(N_281));
    NOR2B \crc_out_ff_RNO[7]  (.A(N_245), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_out_ff_RNO[7]_net_1 ));
    MX2 \crc_init_ff_RNO_0[8]  (.A(\crc_init_ff_3[8] ), .B(
        crc_init_out[8]), .S(un1_crc_init_en_1_0_net_1), .Y(N_139));
    DFN1 \crc_poly_ff[31]  (.D(\crc_poly_ff_RNO[31]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[31]));
    DFN1 crc_init_sel_ff (.D(crc_init_sel_ff_RNI2BI2B_net_1), .CLK(
        FAB_CLK), .Q(crc_init_sel_ff_net_1));
    DFN1 \crc_init_ff[9]  (.D(\crc_init_ff_RNO[9]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_init_out[9]));
    DFN1 \crc_poly_ff[29]  (.D(\crc_poly_ff_RNO[29]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[29]));
    DFN1 \crc_out_ff[4]  (.D(\crc_out_ff_RNO[4]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_out_ff[4]_net_1 ));
    OR2A \crc_init_ff_RNO[15]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_146), .Y(\crc_init_ff_RNO[15]_net_1 ));
    MX2 \crc_init_ff_RNO_0[2]  (.A(\crc_init_ff_3[2] ), .B(
        crc_init_out[2]), .S(un1_crc_init_en_1_0_net_1), .Y(N_133));
    MX2 \crc_init_ff_RNO_0[29]  (.A(\crc_init_ff_3[29] ), .B(
        crc_init_out[29]), .S(un1_crc_init_en_1_net_1), .Y(N_160));
    NOR2B \crc_idr_ff_RNO[5]  (.A(N_235), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_idr_ff_RNO[5]_net_1 ));
    OR2A \crc_poly_ff_RNO[11]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_209), .Y(\crc_poly_ff_RNO[11]_net_1 ));
    MX2 \byte_ff_RNIQIIL[4]  (.A(\byte_ff[4]_net_1 ), .B(
        \buffer_ff[4]_net_1 ), .S(bypass_byte0), .Y(\crc_data_in0[4] ));
    MX2 \crc_out_ff_RNO_0[10]  (.A(\crc_unit_out[10] ), .B(
        \crc_out_ff[10]_net_1 ), .S(state_byte_0[4]), .Y(N_248));
    NOR2B \crc_poly_ff_RNO[19]  (.A(N_217), .B(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .Y(\crc_poly_ff_RNO[19]_net_1 ));
    DFN1 \buffer_ff[2]  (.D(\buffer_ff_RNO[2]_net_1 ), .CLK(FAB_CLK), 
        .Q(\buffer_ff[2]_net_1 ));
    DFN1 \crc_out_ff[7]  (.D(\crc_out_ff_RNO[7]_net_1 ), .CLK(FAB_CLK), 
        .Q(\crc_out_ff[7]_net_1 ));
    OR2A \crc_init_ff_RNO[21]  (.A(crc_ahb_ip_MSS_0_M2F_RESET_N), .B(
        N_152), .Y(\crc_init_ff_RNO[21]_net_1 ));
    DFN1 \crc_poly_ff[1]  (.D(\crc_poly_ff_RNO[1]_net_1 ), .CLK(
        FAB_CLK), .Q(crc_poly_out[1]));
    
endmodule


module crc_unit(
       crc_poly_size,
       state_byte,
       bus_size,
       bus_wr_0,
       bus_wr_1,
       bus_wr_16,
       bus_wr_25,
       bus_wr_2,
       bus_wr_3,
       crc_idr_out,
       crc_out,
       crc_init_out,
       crc_poly_out,
       rev_in_type_0,
       rev_in_type,
       FAB_CLK,
       crc_init_en,
       crc_poly_en,
       N_348,
       N_350,
       N_352,
       N_353,
       crc_poly_en_0,
       N_358,
       N_360,
       N_361,
       N_364,
       N_365,
       N_366,
       N_332,
       N_333,
       N_334,
       N_335,
       N_336,
       N_337,
       crc_idr_en,
       N_347,
       rev_out_type_0,
       rev_out_type,
       crc_ahb_ip_MSS_0_M2F_RESET_N,
       crc_init_en_0,
       N_367,
       crc_poly_size_77,
       N_349,
       N_357,
       N_356,
       N_354,
       N_351,
       N_362,
       N_355,
       N_363,
       crc_poly_size_77_0,
       buffer_write_en,
       buffer_full,
       reset_pending,
       reset_chain
    );
input  [1:0] crc_poly_size;
output [4:4] state_byte;
input  [1:0] bus_size;
input  bus_wr_0;
input  bus_wr_1;
input  bus_wr_16;
input  bus_wr_25;
input  bus_wr_2;
input  bus_wr_3;
output [7:0] crc_idr_out;
output [31:0] crc_out;
output [31:0] crc_init_out;
output [31:0] crc_poly_out;
input  [0:0] rev_in_type_0;
input  [1:0] rev_in_type;
input  FAB_CLK;
input  crc_init_en;
input  crc_poly_en;
input  N_348;
input  N_350;
input  N_352;
input  N_353;
input  crc_poly_en_0;
input  N_358;
input  N_360;
input  N_361;
input  N_364;
input  N_365;
input  N_366;
input  N_332;
input  N_333;
input  N_334;
input  N_335;
input  N_336;
input  N_337;
input  crc_idr_en;
input  N_347;
input  rev_out_type_0;
input  rev_out_type;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;
input  crc_init_en_0;
input  N_367;
output crc_poly_size_77;
input  N_349;
input  N_357;
input  N_356;
input  N_354;
input  N_351;
input  N_362;
input  N_355;
input  N_363;
input  crc_poly_size_77_0;
input  buffer_write_en;
output buffer_full;
output reset_pending;
input  reset_chain;

    wire \state_byte_i[0] , \state_byte_0[4] , \size_in[0] , 
        \size_in[1] , N_56, byte_en_0, byte_en, buffer_en_0, buffer_en, 
        N_118_1, N_128, N_294, bypass_byte0, GND, VCC;
    
    crc_control_unit CONTROL_UNIT (.state_byte_0({\state_byte_0[4] }), 
        .size_in({\size_in[1] , \size_in[0] }), .state_byte_3(
        state_byte[4]), .state_byte_i({\state_byte_i[0] }), .FAB_CLK(
        FAB_CLK), .byte_en_0(byte_en_0), .buffer_en_0(buffer_en_0), 
        .buffer_write_en(buffer_write_en), .buffer_full(buffer_full), 
        .reset_pending(reset_pending), .reset_chain(reset_chain), 
        .N_294(N_294), .crc_ahb_ip_MSS_0_M2F_RESET_N(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .N_128(N_128), .byte_en(byte_en)
        , .N_56(N_56), .bypass_byte0(bypass_byte0), .buffer_en(
        buffer_en), .N_118_1(N_118_1));
    VCC VCC_i (.Y(VCC));
    crc_datapath DATAPATH (.crc_poly_size({crc_poly_size[1], 
        crc_poly_size[0]}), .state_byte_i({\state_byte_i[0] }), 
        .state_byte({state_byte[4]}), .state_byte_0({\state_byte_0[4] })
        , .size_in({\size_in[1] , \size_in[0] }), .bus_size({
        bus_size[1], bus_size[0]}), .bus_wr_0(bus_wr_0), .bus_wr_1(
        bus_wr_1), .bus_wr_16(bus_wr_16), .bus_wr_25(bus_wr_25), 
        .bus_wr_2(bus_wr_2), .bus_wr_3(bus_wr_3), .crc_idr_out({
        crc_idr_out[7], crc_idr_out[6], crc_idr_out[5], crc_idr_out[4], 
        crc_idr_out[3], crc_idr_out[2], crc_idr_out[1], crc_idr_out[0]})
        , .crc_out({crc_out[31], crc_out[30], crc_out[29], crc_out[28], 
        crc_out[27], crc_out[26], crc_out[25], crc_out[24], 
        crc_out[23], crc_out[22], crc_out[21], crc_out[20], 
        crc_out[19], crc_out[18], crc_out[17], crc_out[16], 
        crc_out[15], crc_out[14], crc_out[13], crc_out[12], 
        crc_out[11], crc_out[10], crc_out[9], crc_out[8], crc_out[7], 
        crc_out[6], crc_out[5], crc_out[4], crc_out[3], crc_out[2], 
        crc_out[1], crc_out[0]}), .crc_init_out({crc_init_out[31], 
        crc_init_out[30], crc_init_out[29], crc_init_out[28], 
        crc_init_out[27], crc_init_out[26], crc_init_out[25], 
        crc_init_out[24], crc_init_out[23], crc_init_out[22], 
        crc_init_out[21], crc_init_out[20], crc_init_out[19], 
        crc_init_out[18], crc_init_out[17], crc_init_out[16], 
        crc_init_out[15], crc_init_out[14], crc_init_out[13], 
        crc_init_out[12], crc_init_out[11], crc_init_out[10], 
        crc_init_out[9], crc_init_out[8], crc_init_out[7], 
        crc_init_out[6], crc_init_out[5], crc_init_out[4], 
        crc_init_out[3], crc_init_out[2], crc_init_out[1], 
        crc_init_out[0]}), .crc_poly_out({crc_poly_out[31], 
        crc_poly_out[30], crc_poly_out[29], crc_poly_out[28], 
        crc_poly_out[27], crc_poly_out[26], crc_poly_out[25], 
        crc_poly_out[24], crc_poly_out[23], crc_poly_out[22], 
        crc_poly_out[21], crc_poly_out[20], crc_poly_out[19], 
        crc_poly_out[18], crc_poly_out[17], crc_poly_out[16], 
        crc_poly_out[15], crc_poly_out[14], crc_poly_out[13], 
        crc_poly_out[12], crc_poly_out[11], crc_poly_out[10], 
        crc_poly_out[9], crc_poly_out[8], crc_poly_out[7], 
        crc_poly_out[6], crc_poly_out[5], crc_poly_out[4], 
        crc_poly_out[3], crc_poly_out[2], crc_poly_out[1], 
        crc_poly_out[0]}), .rev_in_type_0({rev_in_type_0[0]}), 
        .rev_in_type({rev_in_type[1], rev_in_type[0]}), .FAB_CLK(
        FAB_CLK), .N_56(N_56), .crc_init_en(crc_init_en), .byte_en_0(
        byte_en_0), .byte_en(byte_en), .crc_poly_en(crc_poly_en), 
        .N_348(N_348), .N_350(N_350), .N_352(N_352), .N_353(N_353), 
        .crc_poly_en_0(crc_poly_en_0), .N_358(N_358), .N_360(N_360), 
        .N_361(N_361), .N_364(N_364), .N_365(N_365), .N_366(N_366), 
        .N_332(N_332), .N_333(N_333), .N_334(N_334), .N_335(N_335), 
        .N_336(N_336), .N_337(N_337), .crc_idr_en(crc_idr_en), .N_347(
        N_347), .buffer_en_0(buffer_en_0), .buffer_en(buffer_en), 
        .rev_out_type_0(rev_out_type_0), .rev_out_type(rev_out_type), 
        .N_118_1(N_118_1), .crc_ahb_ip_MSS_0_M2F_RESET_N(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .N_128(N_128), .N_294_0(N_294), 
        .bypass_byte0(bypass_byte0), .crc_init_en_0(crc_init_en_0), 
        .N_367(N_367), .crc_poly_size_77(crc_poly_size_77), .N_349(
        N_349), .N_357(N_357), .N_356(N_356), .N_354(N_354), .N_351(
        N_351), .N_362(N_362), .N_355(N_355), .N_363(N_363), 
        .crc_poly_size_77_0(crc_poly_size_77_0));
    GND GND_i (.Y(GND));
    
endmodule


module crc_ip(
       HRDATA_2,
       HRDATA_1,
       HRDATA_0_20,
       HRDATA_0_15,
       HRDATA_0_31,
       HRDATA_0_2,
       HRDATA_0_17,
       HRDATA_0_0,
       HRDATA_0_28,
       HRDATA_0_29,
       HRDATA_0_26,
       HRDATA_0_11,
       HRDATA_0_12,
       HRDATA_0_16,
       HRDATA_0_30,
       HRDATA_0_14,
       HRDATA_0_19,
       HRDATA_0_13,
       HRDATA_0_27,
       HRDATA_0_25,
       HRDATA_0_24,
       HRDATA_0_8,
       HRDATA_0_9,
       HRDATA_0_10,
       HRDATA_0_1,
       HRDATA_0_18,
       HRDATA_0_21,
       HRDATA_0_22,
       HRDATA_0_23,
       un4_HRDATA,
       bus_wr_0,
       bus_wr_3,
       bus_wr_1,
       bus_wr_16,
       bus_wr_25,
       bus_wr_2,
       FAB_CLK,
       CoreAHBLite_0_AHBmslave5_HREADY_i_0,
       N_347,
       crc_ahb_ip_MSS_0_M2F_RESET_N,
       N_350,
       N_348,
       N_349,
       un1_masterAddrInProg_6,
       N_5,
       N_408,
       N_409,
       N_387,
       N_340,
       N_341,
       N_342,
       N_352,
       N_353,
       N_358,
       N_360,
       N_361,
       N_364,
       N_365,
       N_366,
       N_332,
       N_333,
       N_334,
       N_335,
       N_336,
       N_337,
       N_367,
       crc_poly_size_77,
       N_357,
       N_356,
       N_354,
       N_351,
       N_362,
       N_355,
       N_363,
       crc_poly_size_77_0
    );
output [7:3] HRDATA_2;
output [7:0] HRDATA_1;
output HRDATA_0_20;
output HRDATA_0_15;
output HRDATA_0_31;
output HRDATA_0_2;
output HRDATA_0_17;
output HRDATA_0_0;
output HRDATA_0_28;
output HRDATA_0_29;
output HRDATA_0_26;
output HRDATA_0_11;
output HRDATA_0_12;
output HRDATA_0_16;
output HRDATA_0_30;
output HRDATA_0_14;
output HRDATA_0_19;
output HRDATA_0_13;
output HRDATA_0_27;
output HRDATA_0_25;
output HRDATA_0_24;
output HRDATA_0_8;
output HRDATA_0_9;
output HRDATA_0_10;
output HRDATA_0_1;
output HRDATA_0_18;
output HRDATA_0_21;
output HRDATA_0_22;
output HRDATA_0_23;
output [31:8] un4_HRDATA;
input  bus_wr_0;
input  bus_wr_3;
input  bus_wr_1;
input  bus_wr_16;
input  bus_wr_25;
input  bus_wr_2;
input  FAB_CLK;
output CoreAHBLite_0_AHBmslave5_HREADY_i_0;
input  N_347;
input  crc_ahb_ip_MSS_0_M2F_RESET_N;
input  N_350;
input  N_348;
input  N_349;
input  un1_masterAddrInProg_6;
input  N_5;
input  N_408;
input  N_409;
input  N_387;
input  N_340;
input  N_341;
input  N_342;
input  N_352;
input  N_353;
input  N_358;
input  N_360;
input  N_361;
input  N_364;
input  N_365;
input  N_366;
input  N_332;
input  N_333;
input  N_334;
input  N_335;
input  N_336;
input  N_337;
input  N_367;
output crc_poly_size_77;
input  N_357;
input  N_356;
input  N_354;
input  N_351;
input  N_362;
input  N_355;
input  N_363;
input  crc_poly_size_77_0;

    wire \rev_in_type_0[0] , \crc_idr_out[0] , \crc_idr_out[1] , 
        \crc_idr_out[2] , \crc_idr_out[3] , \crc_idr_out[4] , 
        \crc_idr_out[5] , \crc_idr_out[6] , \crc_idr_out[7] , 
        \state_byte[4] , \crc_poly_size[0] , \crc_poly_size[1] , 
        \rev_in_type[0] , \rev_in_type[1] , \crc_out[0] , \crc_out[1] , 
        \crc_out[2] , \crc_out[3] , \crc_out[4] , \crc_out[5] , 
        \crc_out[6] , \crc_out[7] , \crc_out[8] , \crc_out[9] , 
        \crc_out[10] , \crc_out[11] , \crc_out[12] , \crc_out[13] , 
        \crc_out[14] , \crc_out[15] , \crc_out[16] , \crc_out[17] , 
        \crc_out[18] , \crc_out[19] , \crc_out[20] , \crc_out[21] , 
        \crc_out[22] , \crc_out[23] , \crc_out[24] , \crc_out[25] , 
        \crc_out[26] , \crc_out[27] , \crc_out[28] , \crc_out[29] , 
        \crc_out[30] , \crc_out[31] , \crc_poly_out[0] , 
        \crc_poly_out[1] , \crc_poly_out[2] , \crc_poly_out[3] , 
        \crc_poly_out[4] , \crc_poly_out[5] , \crc_poly_out[6] , 
        \crc_poly_out[7] , \crc_poly_out[8] , \crc_poly_out[9] , 
        \crc_poly_out[10] , \crc_poly_out[11] , \crc_poly_out[12] , 
        \crc_poly_out[13] , \crc_poly_out[14] , \crc_poly_out[15] , 
        \crc_poly_out[16] , \crc_poly_out[17] , \crc_poly_out[18] , 
        \crc_poly_out[19] , \crc_poly_out[20] , \crc_poly_out[21] , 
        \crc_poly_out[22] , \crc_poly_out[23] , \crc_poly_out[24] , 
        \crc_poly_out[25] , \crc_poly_out[26] , \crc_poly_out[27] , 
        \crc_poly_out[28] , \crc_poly_out[29] , \crc_poly_out[30] , 
        \crc_poly_out[31] , \crc_init_out[0] , \crc_init_out[1] , 
        \crc_init_out[2] , \crc_init_out[3] , \crc_init_out[4] , 
        \crc_init_out[5] , \crc_init_out[6] , \crc_init_out[7] , 
        \crc_init_out[8] , \crc_init_out[9] , \crc_init_out[10] , 
        \crc_init_out[11] , \crc_init_out[12] , \crc_init_out[13] , 
        \crc_init_out[14] , \crc_init_out[15] , \crc_init_out[16] , 
        \crc_init_out[17] , \crc_init_out[18] , \crc_init_out[19] , 
        \crc_init_out[20] , \crc_init_out[21] , \crc_init_out[22] , 
        \crc_init_out[23] , \crc_init_out[24] , \crc_init_out[25] , 
        \crc_init_out[26] , \crc_init_out[27] , \crc_init_out[28] , 
        \crc_init_out[29] , \crc_init_out[30] , \crc_init_out[31] , 
        \bus_size[0] , \bus_size[1] , rev_out_type_0, crc_poly_en_0, 
        crc_init_en_0, buffer_full, buffer_write_en, reset_pending, 
        rev_out_type, reset_chain, crc_poly_en, crc_init_en, 
        crc_idr_en, GND, VCC;
    
    host_interface HOST_INTERFACE (.rev_in_type_0({\rev_in_type_0[0] })
        , .HRDATA_2({HRDATA_2[7], HRDATA_2[6], HRDATA_2[5], 
        HRDATA_2[4], HRDATA_2[3]}), .HRDATA_1({HRDATA_1[7], 
        HRDATA_1[6], HRDATA_1[5], HRDATA_1[4], HRDATA_1[3], 
        HRDATA_1[2], HRDATA_1[1], HRDATA_1[0]}), .crc_idr_out({
        \crc_idr_out[7] , \crc_idr_out[6] , \crc_idr_out[5] , 
        \crc_idr_out[4] , \crc_idr_out[3] , \crc_idr_out[2] , 
        \crc_idr_out[1] , \crc_idr_out[0] }), .HRDATA_0_20(HRDATA_0_20)
        , .HRDATA_0_15(HRDATA_0_15), .HRDATA_0_31(HRDATA_0_31), 
        .HRDATA_0_2(HRDATA_0_2), .HRDATA_0_17(HRDATA_0_17), 
        .HRDATA_0_0(HRDATA_0_0), .HRDATA_0_28(HRDATA_0_28), 
        .HRDATA_0_29(HRDATA_0_29), .HRDATA_0_26(HRDATA_0_26), 
        .HRDATA_0_11(HRDATA_0_11), .HRDATA_0_12(HRDATA_0_12), 
        .HRDATA_0_16(HRDATA_0_16), .HRDATA_0_30(HRDATA_0_30), 
        .HRDATA_0_14(HRDATA_0_14), .HRDATA_0_19(HRDATA_0_19), 
        .HRDATA_0_13(HRDATA_0_13), .HRDATA_0_27(HRDATA_0_27), 
        .HRDATA_0_25(HRDATA_0_25), .HRDATA_0_24(HRDATA_0_24), 
        .HRDATA_0_8(HRDATA_0_8), .HRDATA_0_9(HRDATA_0_9), .HRDATA_0_10(
        HRDATA_0_10), .HRDATA_0_1(HRDATA_0_1), .HRDATA_0_18(
        HRDATA_0_18), .HRDATA_0_21(HRDATA_0_21), .HRDATA_0_22(
        HRDATA_0_22), .HRDATA_0_23(HRDATA_0_23), .state_byte({
        \state_byte[4] }), .crc_poly_size({\crc_poly_size[1] , 
        \crc_poly_size[0] }), .rev_in_type({\rev_in_type[1] , 
        \rev_in_type[0] }), .bus_wr_0(bus_wr_0), .bus_wr_3(bus_wr_3), 
        .crc_out({\crc_out[31] , \crc_out[30] , \crc_out[29] , 
        \crc_out[28] , \crc_out[27] , \crc_out[26] , \crc_out[25] , 
        \crc_out[24] , \crc_out[23] , \crc_out[22] , \crc_out[21] , 
        \crc_out[20] , \crc_out[19] , \crc_out[18] , \crc_out[17] , 
        \crc_out[16] , \crc_out[15] , \crc_out[14] , \crc_out[13] , 
        \crc_out[12] , \crc_out[11] , \crc_out[10] , \crc_out[9] , 
        \crc_out[8] , \crc_out[7] , \crc_out[6] , \crc_out[5] , 
        \crc_out[4] , \crc_out[3] , \crc_out[2] , \crc_out[1] , 
        \crc_out[0] }), .crc_poly_out({\crc_poly_out[31] , 
        \crc_poly_out[30] , \crc_poly_out[29] , \crc_poly_out[28] , 
        \crc_poly_out[27] , \crc_poly_out[26] , \crc_poly_out[25] , 
        \crc_poly_out[24] , \crc_poly_out[23] , \crc_poly_out[22] , 
        \crc_poly_out[21] , \crc_poly_out[20] , \crc_poly_out[19] , 
        \crc_poly_out[18] , \crc_poly_out[17] , \crc_poly_out[16] , 
        \crc_poly_out[15] , \crc_poly_out[14] , \crc_poly_out[13] , 
        \crc_poly_out[12] , \crc_poly_out[11] , \crc_poly_out[10] , 
        \crc_poly_out[9] , \crc_poly_out[8] , \crc_poly_out[7] , 
        \crc_poly_out[6] , \crc_poly_out[5] , \crc_poly_out[4] , 
        \crc_poly_out[3] , \crc_poly_out[2] , \crc_poly_out[1] , 
        \crc_poly_out[0] }), .un4_HRDATA_9(un4_HRDATA[9]), 
        .un4_HRDATA_10(un4_HRDATA[10]), .un4_HRDATA_15(un4_HRDATA[15]), 
        .un4_HRDATA_16(un4_HRDATA[16]), .un4_HRDATA_17(un4_HRDATA[17]), 
        .un4_HRDATA_18(un4_HRDATA[18]), .un4_HRDATA_21(un4_HRDATA[21]), 
        .un4_HRDATA_22(un4_HRDATA[22]), .un4_HRDATA_23(un4_HRDATA[23]), 
        .un4_HRDATA_26(un4_HRDATA[26]), .un4_HRDATA_27(un4_HRDATA[27]), 
        .un4_HRDATA_28(un4_HRDATA[28]), .un4_HRDATA_29(un4_HRDATA[29]), 
        .un4_HRDATA_30(un4_HRDATA[30]), .un4_HRDATA_31(un4_HRDATA[31]), 
        .un4_HRDATA_14(un4_HRDATA[14]), .un4_HRDATA_13(un4_HRDATA[13]), 
        .un4_HRDATA_12(un4_HRDATA[12]), .un4_HRDATA_11(un4_HRDATA[11]), 
        .un4_HRDATA_24(un4_HRDATA[24]), .un4_HRDATA_8(un4_HRDATA[8]), 
        .un4_HRDATA_25(un4_HRDATA[25]), .un4_HRDATA_19(un4_HRDATA[19]), 
        .un4_HRDATA_20(un4_HRDATA[20]), .crc_init_out({
        \crc_init_out[31] , \crc_init_out[30] , \crc_init_out[29] , 
        \crc_init_out[28] , \crc_init_out[27] , \crc_init_out[26] , 
        \crc_init_out[25] , \crc_init_out[24] , \crc_init_out[23] , 
        \crc_init_out[22] , \crc_init_out[21] , \crc_init_out[20] , 
        \crc_init_out[19] , \crc_init_out[18] , \crc_init_out[17] , 
        \crc_init_out[16] , \crc_init_out[15] , \crc_init_out[14] , 
        \crc_init_out[13] , \crc_init_out[12] , \crc_init_out[11] , 
        \crc_init_out[10] , \crc_init_out[9] , \crc_init_out[8] , 
        \crc_init_out[7] , \crc_init_out[6] , \crc_init_out[5] , 
        \crc_init_out[4] , \crc_init_out[3] , \crc_init_out[2] , 
        \crc_init_out[1] , \crc_init_out[0] }), .bus_size({
        \bus_size[1] , \bus_size[0] }), .FAB_CLK(FAB_CLK), 
        .rev_out_type_0(rev_out_type_0), .crc_poly_en_0(crc_poly_en_0), 
        .crc_init_en_0(crc_init_en_0), 
        .CoreAHBLite_0_AHBmslave5_HREADY_i_0(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .N_347(N_347), 
        .buffer_full(buffer_full), .buffer_write_en(buffer_write_en), 
        .reset_pending(reset_pending), .crc_ahb_ip_MSS_0_M2F_RESET_N(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .rev_out_type(rev_out_type), 
        .N_350(N_350), .reset_chain(reset_chain), .crc_poly_en(
        crc_poly_en), .crc_init_en(crc_init_en), .N_348(N_348), .N_349(
        N_349), .crc_idr_en(crc_idr_en), .un1_masterAddrInProg_6(
        un1_masterAddrInProg_6), .N_5(N_5), .N_408(N_408), .N_409(
        N_409), .N_387(N_387), .N_340(N_340), .N_341(N_341), .N_342(
        N_342));
    crc_unit CRC_UNIT (.crc_poly_size({\crc_poly_size[1] , 
        \crc_poly_size[0] }), .state_byte({\state_byte[4] }), 
        .bus_size({\bus_size[1] , \bus_size[0] }), .bus_wr_0(bus_wr_0), 
        .bus_wr_1(bus_wr_1), .bus_wr_16(bus_wr_16), .bus_wr_25(
        bus_wr_25), .bus_wr_2(bus_wr_2), .bus_wr_3(bus_wr_3), 
        .crc_idr_out({\crc_idr_out[7] , \crc_idr_out[6] , 
        \crc_idr_out[5] , \crc_idr_out[4] , \crc_idr_out[3] , 
        \crc_idr_out[2] , \crc_idr_out[1] , \crc_idr_out[0] }), 
        .crc_out({\crc_out[31] , \crc_out[30] , \crc_out[29] , 
        \crc_out[28] , \crc_out[27] , \crc_out[26] , \crc_out[25] , 
        \crc_out[24] , \crc_out[23] , \crc_out[22] , \crc_out[21] , 
        \crc_out[20] , \crc_out[19] , \crc_out[18] , \crc_out[17] , 
        \crc_out[16] , \crc_out[15] , \crc_out[14] , \crc_out[13] , 
        \crc_out[12] , \crc_out[11] , \crc_out[10] , \crc_out[9] , 
        \crc_out[8] , \crc_out[7] , \crc_out[6] , \crc_out[5] , 
        \crc_out[4] , \crc_out[3] , \crc_out[2] , \crc_out[1] , 
        \crc_out[0] }), .crc_init_out({\crc_init_out[31] , 
        \crc_init_out[30] , \crc_init_out[29] , \crc_init_out[28] , 
        \crc_init_out[27] , \crc_init_out[26] , \crc_init_out[25] , 
        \crc_init_out[24] , \crc_init_out[23] , \crc_init_out[22] , 
        \crc_init_out[21] , \crc_init_out[20] , \crc_init_out[19] , 
        \crc_init_out[18] , \crc_init_out[17] , \crc_init_out[16] , 
        \crc_init_out[15] , \crc_init_out[14] , \crc_init_out[13] , 
        \crc_init_out[12] , \crc_init_out[11] , \crc_init_out[10] , 
        \crc_init_out[9] , \crc_init_out[8] , \crc_init_out[7] , 
        \crc_init_out[6] , \crc_init_out[5] , \crc_init_out[4] , 
        \crc_init_out[3] , \crc_init_out[2] , \crc_init_out[1] , 
        \crc_init_out[0] }), .crc_poly_out({\crc_poly_out[31] , 
        \crc_poly_out[30] , \crc_poly_out[29] , \crc_poly_out[28] , 
        \crc_poly_out[27] , \crc_poly_out[26] , \crc_poly_out[25] , 
        \crc_poly_out[24] , \crc_poly_out[23] , \crc_poly_out[22] , 
        \crc_poly_out[21] , \crc_poly_out[20] , \crc_poly_out[19] , 
        \crc_poly_out[18] , \crc_poly_out[17] , \crc_poly_out[16] , 
        \crc_poly_out[15] , \crc_poly_out[14] , \crc_poly_out[13] , 
        \crc_poly_out[12] , \crc_poly_out[11] , \crc_poly_out[10] , 
        \crc_poly_out[9] , \crc_poly_out[8] , \crc_poly_out[7] , 
        \crc_poly_out[6] , \crc_poly_out[5] , \crc_poly_out[4] , 
        \crc_poly_out[3] , \crc_poly_out[2] , \crc_poly_out[1] , 
        \crc_poly_out[0] }), .rev_in_type_0({\rev_in_type_0[0] }), 
        .rev_in_type({\rev_in_type[1] , \rev_in_type[0] }), .FAB_CLK(
        FAB_CLK), .crc_init_en(crc_init_en), .crc_poly_en(crc_poly_en), 
        .N_348(N_348), .N_350(N_350), .N_352(N_352), .N_353(N_353), 
        .crc_poly_en_0(crc_poly_en_0), .N_358(N_358), .N_360(N_360), 
        .N_361(N_361), .N_364(N_364), .N_365(N_365), .N_366(N_366), 
        .N_332(N_332), .N_333(N_333), .N_334(N_334), .N_335(N_335), 
        .N_336(N_336), .N_337(N_337), .crc_idr_en(crc_idr_en), .N_347(
        N_347), .rev_out_type_0(rev_out_type_0), .rev_out_type(
        rev_out_type), .crc_ahb_ip_MSS_0_M2F_RESET_N(
        crc_ahb_ip_MSS_0_M2F_RESET_N), .crc_init_en_0(crc_init_en_0), 
        .N_367(N_367), .crc_poly_size_77(crc_poly_size_77), .N_349(
        N_349), .N_357(N_357), .N_356(N_356), .N_354(N_354), .N_351(
        N_351), .N_362(N_362), .N_355(N_355), .N_363(N_363), 
        .crc_poly_size_77_0(crc_poly_size_77_0), .buffer_write_en(
        buffer_write_en), .buffer_full(buffer_full), .reset_pending(
        reset_pending), .reset_chain(reset_chain));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    
endmodule


module crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC(
       FAB_CLK,
       GLA0
    );
output FAB_CLK;
output GLA0;

    wire N_CLKA_RCOSC, I_MSSCCC_GLA, I_MSSCCC_GLC, I_MSSCCC_LOCK, 
        I_MSSCCC_LOCKMSS, I_MSSCCC_MACCLK, I_MSSCCC_YB, I_MSSCCC_YC, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND;
    
    MSS_CCC #( .VCOFREQUENCY(-1.000000) )  I_MSSCCC (.CLKA(
        N_CLKA_RCOSC), .EXTFB(crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND)
        , .GLA(I_MSSCCC_GLA), .GLAMSS(GLA0), .LOCK(I_MSSCCC_LOCK), 
        .LOCKMSS(I_MSSCCC_LOCKMSS), .CLKB(
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND), .GLB(FAB_CLK), .YB(
        I_MSSCCC_YB), .CLKC(crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND), 
        .GLC(I_MSSCCC_GLC), .YC(I_MSSCCC_YC), .MACCLK(I_MSSCCC_MACCLK), 
        .OADIV({crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .OADIVHALF(
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND), .OAMUX({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .BYPASSA(
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC), .DLYGLA({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .DLYGLAMSS({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .DLYGLAFAB({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .OBDIV({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC}), .OBDIVHALF(
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND), .OBMUX({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC}), .BYPASSB(
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND), .DLYGLB({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .OCDIV({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC}), .OCDIVHALF(
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND), .OCMUX({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .BYPASSC(
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC), .DLYGLC({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .FINDIV({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .FBDIV({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .FBDLY({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC}), .FBSEL({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC}), .XDLYSEL(
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND), .GLMUXSEL({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}), .GLMUXCFG({
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND, 
        crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND}));
    VCC VCC_i (.Y(crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_VCC));
    RCOSC I_RCOSC (.CLKOUT(N_CLKA_RCOSC));
    GND GND_i (.Y(crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC_GND));
    
endmodule


module crc_ahb_ip_MSS(
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_3,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_4,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_18,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_19,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE,
       crc_ahb_ip_MSS_0_M2F_RESET_N,
       defSlaveSMCurrentState_RNI5UNRI,
       UART_0_TXD,
       UART_0_RXD,
       MSS_RESET_N,
       FAB_CLK,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK,
       crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE,
       N_153
    );
output [1:1] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS;
output crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2;
output crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_3;
output crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_4;
output crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16;
output crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17;
output crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_18;
output crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_19;
output [31:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA;
input  [31:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA;
output [1:0] crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE;
output crc_ahb_ip_MSS_0_M2F_RESET_N;
input  defSlaveSMCurrentState_RNI5UNRI;
output UART_0_TXD;
input  UART_0_RXD;
input  MSS_RESET_N;
output FAB_CLK;
output crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK;
output crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE;
input  N_153;

    wire MSS_ADLIB_INST_M2FRESETn, N_266, MSS_UART_0_TXD_D, 
        MSS_UART_0_RXD_Y, MSS_RESET_0_MSS_RESET_N_Y, 
        MSS_ADLIB_INST_EMCRWn, MSS_ADLIB_INST_EMCDBOE, 
        MSS_ADLIB_INST_EMCCLK, crc_ahb_ip_MSS_VCC, 
        MSS_ADLIB_INST_CALIBOUT, crc_ahb_ip_MSS_GND, 
        MSS_ADLIB_INST_WDINT, MSS_ADLIB_INST_DEEPSLEEP, 
        MSS_ADLIB_INST_SLEEP, MSS_ADLIB_INST_TXEV, 
        MSS_ADLIB_INST_UART0RTSn, MSS_ADLIB_INST_UART0DTRn, 
        MSS_ADLIB_INST_UART1RTSn, MSS_ADLIB_INST_UART1DTRn, 
        MSS_ADLIB_INST_I2C0SMBUSNO, MSS_ADLIB_INST_I2C1SMBUSNO, 
        MSS_ADLIB_INST_I2C0SMBALERTNO, MSS_ADLIB_INST_I2C1SMBALERTNO, 
        GLA0, MSS_ADLIB_INST_SPI0DO, MSS_ADLIB_INST_SPI0DOE, 
        MSS_ADLIB_INST_SPI0CLKO, MSS_ADLIB_INST_SPI0MODE, 
        MSS_ADLIB_INST_I2C0SDAO, MSS_ADLIB_INST_I2C0SCLO, 
        MSS_ADLIB_INST_SPI1DO, MSS_ADLIB_INST_SPI1DOE, 
        MSS_ADLIB_INST_SPI1CLKO, MSS_ADLIB_INST_SPI1MODE, 
        MSS_ADLIB_INST_UART1TXD, MSS_ADLIB_INST_I2C1SDAO, 
        MSS_ADLIB_INST_I2C1SCLO, MSS_ADLIB_INST_MACTXEN, 
        MSS_ADLIB_INST_MACMDO, MSS_ADLIB_INST_MACMDEN, 
        MSS_ADLIB_INST_MACMDC, \MSS_ADLIB_INST_MACM2FTXD[0] , 
        \MSS_ADLIB_INST_MACM2FTXD[1] , MSS_ADLIB_INST_MACM2FTXEN, 
        MSS_ADLIB_INST_MACM2FMDO, MSS_ADLIB_INST_MACM2FMDEN, 
        MSS_ADLIB_INST_MACM2FMDC, MSS_ADLIB_INST_PUFABn, 
        MSS_ADLIB_INST_FABHREADYOUT, \MSSHTRANS[0] , 
        MSS_ADLIB_INST_LVTTL3, MSS_ADLIB_INST_LVTTL6, 
        MSS_ADLIB_INST_VAREFOUT, MSS_ADLIB_INST_LVTTL1, 
        MSS_ADLIB_INST_SDD2, MSS_ADLIB_INST_LVTTL9, 
        MSS_ADLIB_INST_LVTTL2, MSS_ADLIB_INST_SDD1, 
        MSS_ADLIB_INST_LVTTL5, MSS_ADLIB_INST_SDD0, 
        MSS_ADLIB_INST_LVTTL10, MSS_ADLIB_INST_LVTTL8, 
        MSS_ADLIB_INST_LVTTL0, MSS_ADLIB_INST_LVTTL7, 
        MSS_ADLIB_INST_LVTTL4, MSS_ADLIB_INST_LVTTL11, 
        MSS_ADLIB_INST_FABHRESP, MSS_ADLIB_INST_CMP0, 
        MSS_ADLIB_INST_CMP1, MSS_ADLIB_INST_CMP2, MSS_ADLIB_INST_CMP3, 
        MSS_ADLIB_INST_CMP4, MSS_ADLIB_INST_CMP5, MSS_ADLIB_INST_CMP6, 
        MSS_ADLIB_INST_CMP7, MSS_ADLIB_INST_CMP8, MSS_ADLIB_INST_CMP9, 
        MSS_ADLIB_INST_CMP10, MSS_ADLIB_INST_CMP11, 
        MSS_ADLIB_INST_VCC15GOOD, MSS_ADLIB_INST_VCC33GOOD, 
        \MSS_ADLIB_INST_EMCBYTEN[0] , \MSS_ADLIB_INST_EMCBYTEN[1] , 
        \MSS_ADLIB_INST_EMCAB[0] , \MSS_ADLIB_INST_EMCAB[1] , 
        \MSS_ADLIB_INST_EMCAB[2] , \MSS_ADLIB_INST_EMCAB[3] , 
        \MSS_ADLIB_INST_EMCAB[4] , \MSS_ADLIB_INST_EMCAB[5] , 
        \MSS_ADLIB_INST_EMCAB[6] , \MSS_ADLIB_INST_EMCAB[7] , 
        \MSS_ADLIB_INST_EMCAB[8] , \MSS_ADLIB_INST_EMCAB[9] , 
        \MSS_ADLIB_INST_EMCAB[10] , \MSS_ADLIB_INST_EMCAB[11] , 
        \MSS_ADLIB_INST_EMCAB[12] , \MSS_ADLIB_INST_EMCAB[13] , 
        \MSS_ADLIB_INST_EMCAB[14] , \MSS_ADLIB_INST_EMCAB[15] , 
        \MSS_ADLIB_INST_EMCAB[16] , \MSS_ADLIB_INST_EMCAB[17] , 
        \MSS_ADLIB_INST_EMCAB[18] , \MSS_ADLIB_INST_EMCAB[19] , 
        \MSS_ADLIB_INST_EMCAB[20] , \MSS_ADLIB_INST_EMCAB[21] , 
        \MSS_ADLIB_INST_EMCAB[22] , \MSS_ADLIB_INST_EMCAB[23] , 
        \MSS_ADLIB_INST_EMCAB[24] , \MSS_ADLIB_INST_EMCAB[25] , 
        MSS_ADLIB_INST_EMCOEN0n, MSS_ADLIB_INST_EMCOEN1n, 
        \MSS_ADLIB_INST_EMCWDB[0] , \MSS_ADLIB_INST_EMCWDB[1] , 
        \MSS_ADLIB_INST_EMCWDB[2] , \MSS_ADLIB_INST_EMCWDB[3] , 
        \MSS_ADLIB_INST_EMCWDB[4] , \MSS_ADLIB_INST_EMCWDB[5] , 
        \MSS_ADLIB_INST_EMCWDB[6] , \MSS_ADLIB_INST_EMCWDB[7] , 
        \MSS_ADLIB_INST_EMCWDB[8] , \MSS_ADLIB_INST_EMCWDB[9] , 
        \MSS_ADLIB_INST_EMCWDB[10] , \MSS_ADLIB_INST_EMCWDB[11] , 
        \MSS_ADLIB_INST_EMCWDB[12] , \MSS_ADLIB_INST_EMCWDB[13] , 
        \MSS_ADLIB_INST_EMCWDB[14] , \MSS_ADLIB_INST_EMCWDB[15] , 
        MSS_ADLIB_INST_EMCCS0n, MSS_ADLIB_INST_EMCCS1n, 
        \MSS_ADLIB_INST_GPOE[0] , \MSS_ADLIB_INST_GPOE[1] , 
        \MSS_ADLIB_INST_GPOE[2] , \MSS_ADLIB_INST_GPOE[3] , 
        \MSS_ADLIB_INST_GPOE[4] , \MSS_ADLIB_INST_GPOE[5] , 
        \MSS_ADLIB_INST_GPOE[6] , \MSS_ADLIB_INST_GPOE[7] , 
        \MSS_ADLIB_INST_GPOE[8] , \MSS_ADLIB_INST_GPOE[9] , 
        \MSS_ADLIB_INST_GPOE[10] , \MSS_ADLIB_INST_GPOE[11] , 
        \MSS_ADLIB_INST_GPOE[12] , \MSS_ADLIB_INST_GPOE[13] , 
        \MSS_ADLIB_INST_GPOE[14] , \MSS_ADLIB_INST_GPOE[15] , 
        \MSS_ADLIB_INST_GPOE[16] , \MSS_ADLIB_INST_GPOE[17] , 
        \MSS_ADLIB_INST_GPOE[18] , \MSS_ADLIB_INST_GPOE[19] , 
        \MSS_ADLIB_INST_GPOE[20] , \MSS_ADLIB_INST_GPOE[21] , 
        \MSS_ADLIB_INST_GPOE[22] , \MSS_ADLIB_INST_GPOE[23] , 
        \MSS_ADLIB_INST_GPOE[24] , \MSS_ADLIB_INST_GPOE[25] , 
        \MSS_ADLIB_INST_GPOE[26] , \MSS_ADLIB_INST_GPOE[27] , 
        \MSS_ADLIB_INST_GPOE[28] , \MSS_ADLIB_INST_GPOE[29] , 
        \MSS_ADLIB_INST_GPOE[30] , \MSS_ADLIB_INST_GPOE[31] , 
        \MSS_ADLIB_INST_GPO[0] , \MSS_ADLIB_INST_GPO[1] , 
        \MSS_ADLIB_INST_GPO[2] , \MSS_ADLIB_INST_GPO[3] , 
        \MSS_ADLIB_INST_GPO[4] , \MSS_ADLIB_INST_GPO[5] , 
        \MSS_ADLIB_INST_GPO[6] , \MSS_ADLIB_INST_GPO[7] , 
        \MSS_ADLIB_INST_GPO[8] , \MSS_ADLIB_INST_GPO[9] , 
        \MSS_ADLIB_INST_GPO[10] , \MSS_ADLIB_INST_GPO[11] , 
        \MSS_ADLIB_INST_GPO[12] , \MSS_ADLIB_INST_GPO[13] , 
        \MSS_ADLIB_INST_GPO[14] , \MSS_ADLIB_INST_GPO[15] , 
        \MSS_ADLIB_INST_GPO[16] , \MSS_ADLIB_INST_GPO[17] , 
        \MSS_ADLIB_INST_GPO[18] , \MSS_ADLIB_INST_GPO[19] , 
        \MSS_ADLIB_INST_GPO[20] , \MSS_ADLIB_INST_GPO[21] , 
        \MSS_ADLIB_INST_GPO[22] , \MSS_ADLIB_INST_GPO[23] , 
        \MSS_ADLIB_INST_GPO[24] , \MSS_ADLIB_INST_GPO[25] , 
        \MSS_ADLIB_INST_GPO[26] , \MSS_ADLIB_INST_GPO[27] , 
        \MSS_ADLIB_INST_GPO[28] , \MSS_ADLIB_INST_GPO[29] , 
        \MSS_ADLIB_INST_GPO[30] , \MSS_ADLIB_INST_GPO[31] , 
        \MSS_ADLIB_INST_MSSINT[0] , \MSS_ADLIB_INST_MSSINT[1] , 
        \MSS_ADLIB_INST_MSSINT[2] , \MSS_ADLIB_INST_MSSINT[3] , 
        \MSS_ADLIB_INST_MSSINT[4] , \MSS_ADLIB_INST_MSSINT[5] , 
        \MSS_ADLIB_INST_MSSINT[6] , \MSS_ADLIB_INST_MSSINT[7] , 
        \MSS_ADLIB_INST_SPI0SSO[0] , \MSS_ADLIB_INST_SPI0SSO[1] , 
        \MSS_ADLIB_INST_SPI0SSO[2] , \MSS_ADLIB_INST_SPI0SSO[3] , 
        \MSS_ADLIB_INST_SPI0SSO[4] , \MSS_ADLIB_INST_SPI0SSO[5] , 
        \MSS_ADLIB_INST_SPI0SSO[6] , \MSS_ADLIB_INST_SPI0SSO[7] , 
        \MSS_ADLIB_INST_SPI1SSO[0] , \MSS_ADLIB_INST_SPI1SSO[1] , 
        \MSS_ADLIB_INST_SPI1SSO[2] , \MSS_ADLIB_INST_SPI1SSO[3] , 
        \MSS_ADLIB_INST_SPI1SSO[4] , \MSS_ADLIB_INST_SPI1SSO[5] , 
        \MSS_ADLIB_INST_SPI1SSO[6] , \MSS_ADLIB_INST_SPI1SSO[7] , 
        \MSS_ADLIB_INST_MACTXD[0] , \MSS_ADLIB_INST_MACTXD[1] , 
        \MSS_ADLIB_INST_FABHRDATA[0] , \MSS_ADLIB_INST_FABHRDATA[1] , 
        \MSS_ADLIB_INST_FABHRDATA[2] , \MSS_ADLIB_INST_FABHRDATA[3] , 
        \MSS_ADLIB_INST_FABHRDATA[4] , \MSS_ADLIB_INST_FABHRDATA[5] , 
        \MSS_ADLIB_INST_FABHRDATA[6] , \MSS_ADLIB_INST_FABHRDATA[7] , 
        \MSS_ADLIB_INST_FABHRDATA[8] , \MSS_ADLIB_INST_FABHRDATA[9] , 
        \MSS_ADLIB_INST_FABHRDATA[10] , \MSS_ADLIB_INST_FABHRDATA[11] , 
        \MSS_ADLIB_INST_FABHRDATA[12] , \MSS_ADLIB_INST_FABHRDATA[13] , 
        \MSS_ADLIB_INST_FABHRDATA[14] , \MSS_ADLIB_INST_FABHRDATA[15] , 
        \MSS_ADLIB_INST_FABHRDATA[16] , \MSS_ADLIB_INST_FABHRDATA[17] , 
        \MSS_ADLIB_INST_FABHRDATA[18] , \MSS_ADLIB_INST_FABHRDATA[19] , 
        \MSS_ADLIB_INST_FABHRDATA[20] , \MSS_ADLIB_INST_FABHRDATA[21] , 
        \MSS_ADLIB_INST_FABHRDATA[22] , \MSS_ADLIB_INST_FABHRDATA[23] , 
        \MSS_ADLIB_INST_FABHRDATA[24] , \MSS_ADLIB_INST_FABHRDATA[25] , 
        \MSS_ADLIB_INST_FABHRDATA[26] , \MSS_ADLIB_INST_FABHRDATA[27] , 
        \MSS_ADLIB_INST_FABHRDATA[28] , \MSS_ADLIB_INST_FABHRDATA[29] , 
        \MSS_ADLIB_INST_FABHRDATA[30] , \MSS_ADLIB_INST_FABHRDATA[31] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[0] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[5] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[6] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[7] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[8] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[9] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[10] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[11] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[12] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[13] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[14] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[15] , 
        \MSS_ADLIB_INST_ACEFLAGS[0] , \MSS_ADLIB_INST_ACEFLAGS[1] , 
        \MSS_ADLIB_INST_ACEFLAGS[2] , \MSS_ADLIB_INST_ACEFLAGS[3] , 
        \MSS_ADLIB_INST_ACEFLAGS[4] , \MSS_ADLIB_INST_ACEFLAGS[5] , 
        \MSS_ADLIB_INST_ACEFLAGS[6] , \MSS_ADLIB_INST_ACEFLAGS[7] , 
        \MSS_ADLIB_INST_ACEFLAGS[8] , \MSS_ADLIB_INST_ACEFLAGS[9] , 
        \MSS_ADLIB_INST_ACEFLAGS[10] , \MSS_ADLIB_INST_ACEFLAGS[11] , 
        \MSS_ADLIB_INST_ACEFLAGS[12] , \MSS_ADLIB_INST_ACEFLAGS[13] , 
        \MSS_ADLIB_INST_ACEFLAGS[14] , \MSS_ADLIB_INST_ACEFLAGS[15] , 
        \MSS_ADLIB_INST_ACEFLAGS[16] , \MSS_ADLIB_INST_ACEFLAGS[17] , 
        \MSS_ADLIB_INST_ACEFLAGS[18] , \MSS_ADLIB_INST_ACEFLAGS[19] , 
        \MSS_ADLIB_INST_ACEFLAGS[20] , \MSS_ADLIB_INST_ACEFLAGS[21] , 
        \MSS_ADLIB_INST_ACEFLAGS[22] , \MSS_ADLIB_INST_ACEFLAGS[23] , 
        \MSS_ADLIB_INST_ACEFLAGS[24] , \MSS_ADLIB_INST_ACEFLAGS[25] , 
        \MSS_ADLIB_INST_ACEFLAGS[26] , \MSS_ADLIB_INST_ACEFLAGS[27] , 
        \MSS_ADLIB_INST_ACEFLAGS[28] , \MSS_ADLIB_INST_ACEFLAGS[29] , 
        \MSS_ADLIB_INST_ACEFLAGS[30] , \MSS_ADLIB_INST_ACEFLAGS[31] ;
    
    INBUF_MSS #( .ACT_CONFIG(0), .ACT_PIN("R1") )  
        MSS_RESET_0_MSS_RESET_N (.PAD(MSS_RESET_N), .Y(
        MSS_RESET_0_MSS_RESET_N_Y));
    CLKINT MSS_ADLIB_INST_RNIKNK2 (.A(MSS_ADLIB_INST_M2FRESETn), .Y(
        crc_ahb_ip_MSS_0_M2F_RESET_N));
    OUTBUF_MSS #( .ACT_CONFIG(0), .ACT_PIN("Y22") )  MSS_UART_0_TXD (
        .D(MSS_UART_0_TXD_D), .PAD(UART_0_TXD));
    crc_ahb_ip_MSS_tmp_MSS_CCC_0_MSS_CCC MSS_CCC_0 (.FAB_CLK(FAB_CLK), 
        .GLA0(GLA0));
    INV MSS_ADLIB_INST_RNO (.A(defSlaveSMCurrentState_RNI5UNRI), .Y(
        N_266));
    MSS_AHB #( .ACT_CONFIG(256), .ACT_FCLK(100000000), .ACT_DIE("IP4X3M1")
        , .ACT_PKG("fg484") )  MSS_ADLIB_INST (.MSSHADDR({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_19, 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_18, 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17, 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16, 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[15] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[14] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[13] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[12] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[11] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[10] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[9] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[8] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[7] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[6] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[5] , 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_4, 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_3, 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2, 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[0] }), .MSSHWDATA({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[31], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[30], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[29], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[28], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[27], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[26], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[25], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[24], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[23], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[22], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[21], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[20], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[19], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[18], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[17], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[16], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[15], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[14], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[13], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[12], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[11], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[10], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[9], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[8], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[7], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[6], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[5], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[4], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[3], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[2], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[1], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[0]}), .MSSHTRANS({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS[1], \MSSHTRANS[0] })
        , .MSSHSIZE({crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[1], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[0]}), .MSSHLOCK(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK), .MSSHWRITE(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE), .MSSHRDATA({
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[31], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[30], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[29], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[28], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[27], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[26], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[25], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[24], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[23], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[22], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[21], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[20], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[19], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[18], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[17], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[16], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[15], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[14], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[13], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[12], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[11], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[10], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[9], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[8], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[7], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[6], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[5], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[4], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[3], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[2], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[1], 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[0]}), .MSSHREADY(
        N_266), .MSSHRESP(N_153), .FABHADDR({crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND}), .FABHWDATA({crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND}), .FABHTRANS({crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND}), .FABHSIZE({crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND}), .FABHMASTLOCK(crc_ahb_ip_MSS_GND), 
        .FABHWRITE(crc_ahb_ip_MSS_GND), .FABHSEL(crc_ahb_ip_MSS_GND), 
        .FABHREADY(crc_ahb_ip_MSS_VCC), .FABHRDATA({
        \MSS_ADLIB_INST_FABHRDATA[31] , \MSS_ADLIB_INST_FABHRDATA[30] , 
        \MSS_ADLIB_INST_FABHRDATA[29] , \MSS_ADLIB_INST_FABHRDATA[28] , 
        \MSS_ADLIB_INST_FABHRDATA[27] , \MSS_ADLIB_INST_FABHRDATA[26] , 
        \MSS_ADLIB_INST_FABHRDATA[25] , \MSS_ADLIB_INST_FABHRDATA[24] , 
        \MSS_ADLIB_INST_FABHRDATA[23] , \MSS_ADLIB_INST_FABHRDATA[22] , 
        \MSS_ADLIB_INST_FABHRDATA[21] , \MSS_ADLIB_INST_FABHRDATA[20] , 
        \MSS_ADLIB_INST_FABHRDATA[19] , \MSS_ADLIB_INST_FABHRDATA[18] , 
        \MSS_ADLIB_INST_FABHRDATA[17] , \MSS_ADLIB_INST_FABHRDATA[16] , 
        \MSS_ADLIB_INST_FABHRDATA[15] , \MSS_ADLIB_INST_FABHRDATA[14] , 
        \MSS_ADLIB_INST_FABHRDATA[13] , \MSS_ADLIB_INST_FABHRDATA[12] , 
        \MSS_ADLIB_INST_FABHRDATA[11] , \MSS_ADLIB_INST_FABHRDATA[10] , 
        \MSS_ADLIB_INST_FABHRDATA[9] , \MSS_ADLIB_INST_FABHRDATA[8] , 
        \MSS_ADLIB_INST_FABHRDATA[7] , \MSS_ADLIB_INST_FABHRDATA[6] , 
        \MSS_ADLIB_INST_FABHRDATA[5] , \MSS_ADLIB_INST_FABHRDATA[4] , 
        \MSS_ADLIB_INST_FABHRDATA[3] , \MSS_ADLIB_INST_FABHRDATA[2] , 
        \MSS_ADLIB_INST_FABHRDATA[1] , \MSS_ADLIB_INST_FABHRDATA[0] }), 
        .FABHREADYOUT(MSS_ADLIB_INST_FABHREADYOUT), .FABHRESP(
        MSS_ADLIB_INST_FABHRESP), .SYNCCLKFDBK(FAB_CLK), .CALIBOUT(
        MSS_ADLIB_INST_CALIBOUT), .CALIBIN(crc_ahb_ip_MSS_GND), 
        .FABINT(crc_ahb_ip_MSS_GND), .MSSINT({
        \MSS_ADLIB_INST_MSSINT[7] , \MSS_ADLIB_INST_MSSINT[6] , 
        \MSS_ADLIB_INST_MSSINT[5] , \MSS_ADLIB_INST_MSSINT[4] , 
        \MSS_ADLIB_INST_MSSINT[3] , \MSS_ADLIB_INST_MSSINT[2] , 
        \MSS_ADLIB_INST_MSSINT[1] , \MSS_ADLIB_INST_MSSINT[0] }), 
        .WDINT(MSS_ADLIB_INST_WDINT), .F2MRESETn(crc_ahb_ip_MSS_VCC), 
        .DMAREADY({crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND}), .RXEV(
        crc_ahb_ip_MSS_GND), .VRON(crc_ahb_ip_MSS_GND), .M2FRESETn(
        MSS_ADLIB_INST_M2FRESETn), .DEEPSLEEP(MSS_ADLIB_INST_DEEPSLEEP)
        , .SLEEP(MSS_ADLIB_INST_SLEEP), .TXEV(MSS_ADLIB_INST_TXEV), 
        .GPI({crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND}), 
        .GPO({\MSS_ADLIB_INST_GPO[31] , \MSS_ADLIB_INST_GPO[30] , 
        \MSS_ADLIB_INST_GPO[29] , \MSS_ADLIB_INST_GPO[28] , 
        \MSS_ADLIB_INST_GPO[27] , \MSS_ADLIB_INST_GPO[26] , 
        \MSS_ADLIB_INST_GPO[25] , \MSS_ADLIB_INST_GPO[24] , 
        \MSS_ADLIB_INST_GPO[23] , \MSS_ADLIB_INST_GPO[22] , 
        \MSS_ADLIB_INST_GPO[21] , \MSS_ADLIB_INST_GPO[20] , 
        \MSS_ADLIB_INST_GPO[19] , \MSS_ADLIB_INST_GPO[18] , 
        \MSS_ADLIB_INST_GPO[17] , \MSS_ADLIB_INST_GPO[16] , 
        \MSS_ADLIB_INST_GPO[15] , \MSS_ADLIB_INST_GPO[14] , 
        \MSS_ADLIB_INST_GPO[13] , \MSS_ADLIB_INST_GPO[12] , 
        \MSS_ADLIB_INST_GPO[11] , \MSS_ADLIB_INST_GPO[10] , 
        \MSS_ADLIB_INST_GPO[9] , \MSS_ADLIB_INST_GPO[8] , 
        \MSS_ADLIB_INST_GPO[7] , \MSS_ADLIB_INST_GPO[6] , 
        \MSS_ADLIB_INST_GPO[5] , \MSS_ADLIB_INST_GPO[4] , 
        \MSS_ADLIB_INST_GPO[3] , \MSS_ADLIB_INST_GPO[2] , 
        \MSS_ADLIB_INST_GPO[1] , \MSS_ADLIB_INST_GPO[0] }), .UART0CTSn(
        crc_ahb_ip_MSS_GND), .UART0DSRn(crc_ahb_ip_MSS_GND), .UART0RIn(
        crc_ahb_ip_MSS_GND), .UART0DCDn(crc_ahb_ip_MSS_GND), 
        .UART0RTSn(MSS_ADLIB_INST_UART0RTSn), .UART0DTRn(
        MSS_ADLIB_INST_UART0DTRn), .UART1CTSn(crc_ahb_ip_MSS_GND), 
        .UART1DSRn(crc_ahb_ip_MSS_GND), .UART1RIn(crc_ahb_ip_MSS_GND), 
        .UART1DCDn(crc_ahb_ip_MSS_GND), .UART1RTSn(
        MSS_ADLIB_INST_UART1RTSn), .UART1DTRn(MSS_ADLIB_INST_UART1DTRn)
        , .I2C0SMBUSNI(crc_ahb_ip_MSS_GND), .I2C0SMBALERTNI(
        crc_ahb_ip_MSS_GND), .I2C0BCLK(crc_ahb_ip_MSS_GND), 
        .I2C0SMBUSNO(MSS_ADLIB_INST_I2C0SMBUSNO), .I2C0SMBALERTNO(
        MSS_ADLIB_INST_I2C0SMBALERTNO), .I2C1SMBUSNI(
        crc_ahb_ip_MSS_GND), .I2C1SMBALERTNI(crc_ahb_ip_MSS_GND), 
        .I2C1BCLK(crc_ahb_ip_MSS_GND), .I2C1SMBUSNO(
        MSS_ADLIB_INST_I2C1SMBUSNO), .I2C1SMBALERTNO(
        MSS_ADLIB_INST_I2C1SMBALERTNO), .MACM2FTXD({
        \MSS_ADLIB_INST_MACM2FTXD[1] , \MSS_ADLIB_INST_MACM2FTXD[0] }), 
        .MACF2MRXD({crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND}), 
        .MACM2FTXEN(MSS_ADLIB_INST_MACM2FTXEN), .MACF2MCRSDV(
        crc_ahb_ip_MSS_GND), .MACF2MRXER(crc_ahb_ip_MSS_GND), 
        .MACF2MMDI(crc_ahb_ip_MSS_GND), .MACM2FMDO(
        MSS_ADLIB_INST_MACM2FMDO), .MACM2FMDEN(
        MSS_ADLIB_INST_MACM2FMDEN), .MACM2FMDC(
        MSS_ADLIB_INST_MACM2FMDC), .FABSDD0D(crc_ahb_ip_MSS_GND), 
        .FABSDD1D(crc_ahb_ip_MSS_GND), .FABSDD2D(crc_ahb_ip_MSS_GND), 
        .FABSDD0CLK(crc_ahb_ip_MSS_GND), .FABSDD1CLK(
        crc_ahb_ip_MSS_GND), .FABSDD2CLK(crc_ahb_ip_MSS_GND), 
        .FABACETRIG(crc_ahb_ip_MSS_GND), .ACEFLAGS({
        \MSS_ADLIB_INST_ACEFLAGS[31] , \MSS_ADLIB_INST_ACEFLAGS[30] , 
        \MSS_ADLIB_INST_ACEFLAGS[29] , \MSS_ADLIB_INST_ACEFLAGS[28] , 
        \MSS_ADLIB_INST_ACEFLAGS[27] , \MSS_ADLIB_INST_ACEFLAGS[26] , 
        \MSS_ADLIB_INST_ACEFLAGS[25] , \MSS_ADLIB_INST_ACEFLAGS[24] , 
        \MSS_ADLIB_INST_ACEFLAGS[23] , \MSS_ADLIB_INST_ACEFLAGS[22] , 
        \MSS_ADLIB_INST_ACEFLAGS[21] , \MSS_ADLIB_INST_ACEFLAGS[20] , 
        \MSS_ADLIB_INST_ACEFLAGS[19] , \MSS_ADLIB_INST_ACEFLAGS[18] , 
        \MSS_ADLIB_INST_ACEFLAGS[17] , \MSS_ADLIB_INST_ACEFLAGS[16] , 
        \MSS_ADLIB_INST_ACEFLAGS[15] , \MSS_ADLIB_INST_ACEFLAGS[14] , 
        \MSS_ADLIB_INST_ACEFLAGS[13] , \MSS_ADLIB_INST_ACEFLAGS[12] , 
        \MSS_ADLIB_INST_ACEFLAGS[11] , \MSS_ADLIB_INST_ACEFLAGS[10] , 
        \MSS_ADLIB_INST_ACEFLAGS[9] , \MSS_ADLIB_INST_ACEFLAGS[8] , 
        \MSS_ADLIB_INST_ACEFLAGS[7] , \MSS_ADLIB_INST_ACEFLAGS[6] , 
        \MSS_ADLIB_INST_ACEFLAGS[5] , \MSS_ADLIB_INST_ACEFLAGS[4] , 
        \MSS_ADLIB_INST_ACEFLAGS[3] , \MSS_ADLIB_INST_ACEFLAGS[2] , 
        \MSS_ADLIB_INST_ACEFLAGS[1] , \MSS_ADLIB_INST_ACEFLAGS[0] }), 
        .CMP0(MSS_ADLIB_INST_CMP0), .CMP1(MSS_ADLIB_INST_CMP1), .CMP2(
        MSS_ADLIB_INST_CMP2), .CMP3(MSS_ADLIB_INST_CMP3), .CMP4(
        MSS_ADLIB_INST_CMP4), .CMP5(MSS_ADLIB_INST_CMP5), .CMP6(
        MSS_ADLIB_INST_CMP6), .CMP7(MSS_ADLIB_INST_CMP7), .CMP8(
        MSS_ADLIB_INST_CMP8), .CMP9(MSS_ADLIB_INST_CMP9), .CMP10(
        MSS_ADLIB_INST_CMP10), .CMP11(MSS_ADLIB_INST_CMP11), .LVTTL0EN(
        crc_ahb_ip_MSS_GND), .LVTTL1EN(crc_ahb_ip_MSS_GND), .LVTTL2EN(
        crc_ahb_ip_MSS_GND), .LVTTL3EN(crc_ahb_ip_MSS_GND), .LVTTL4EN(
        crc_ahb_ip_MSS_GND), .LVTTL5EN(crc_ahb_ip_MSS_GND), .LVTTL6EN(
        crc_ahb_ip_MSS_GND), .LVTTL7EN(crc_ahb_ip_MSS_GND), .LVTTL8EN(
        crc_ahb_ip_MSS_GND), .LVTTL9EN(crc_ahb_ip_MSS_GND), .LVTTL10EN(
        crc_ahb_ip_MSS_GND), .LVTTL11EN(crc_ahb_ip_MSS_GND), .LVTTL0(
        MSS_ADLIB_INST_LVTTL0), .LVTTL1(MSS_ADLIB_INST_LVTTL1), 
        .LVTTL2(MSS_ADLIB_INST_LVTTL2), .LVTTL3(MSS_ADLIB_INST_LVTTL3), 
        .LVTTL4(MSS_ADLIB_INST_LVTTL4), .LVTTL5(MSS_ADLIB_INST_LVTTL5), 
        .LVTTL6(MSS_ADLIB_INST_LVTTL6), .LVTTL7(MSS_ADLIB_INST_LVTTL7), 
        .LVTTL8(MSS_ADLIB_INST_LVTTL8), .LVTTL9(MSS_ADLIB_INST_LVTTL9), 
        .LVTTL10(MSS_ADLIB_INST_LVTTL10), .LVTTL11(
        MSS_ADLIB_INST_LVTTL11), .PUFABn(MSS_ADLIB_INST_PUFABn), 
        .VCC15GOOD(MSS_ADLIB_INST_VCC15GOOD), .VCC33GOOD(
        MSS_ADLIB_INST_VCC33GOOD), .FCLK(GLA0), .MACCLKCCC(
        crc_ahb_ip_MSS_GND), .RCOSC(crc_ahb_ip_MSS_GND), .MACCLK(
        crc_ahb_ip_MSS_GND), .PLLLOCK(crc_ahb_ip_MSS_GND), .MSSRESETn(
        MSS_RESET_0_MSS_RESET_N_Y), .GPOE({\MSS_ADLIB_INST_GPOE[31] , 
        \MSS_ADLIB_INST_GPOE[30] , \MSS_ADLIB_INST_GPOE[29] , 
        \MSS_ADLIB_INST_GPOE[28] , \MSS_ADLIB_INST_GPOE[27] , 
        \MSS_ADLIB_INST_GPOE[26] , \MSS_ADLIB_INST_GPOE[25] , 
        \MSS_ADLIB_INST_GPOE[24] , \MSS_ADLIB_INST_GPOE[23] , 
        \MSS_ADLIB_INST_GPOE[22] , \MSS_ADLIB_INST_GPOE[21] , 
        \MSS_ADLIB_INST_GPOE[20] , \MSS_ADLIB_INST_GPOE[19] , 
        \MSS_ADLIB_INST_GPOE[18] , \MSS_ADLIB_INST_GPOE[17] , 
        \MSS_ADLIB_INST_GPOE[16] , \MSS_ADLIB_INST_GPOE[15] , 
        \MSS_ADLIB_INST_GPOE[14] , \MSS_ADLIB_INST_GPOE[13] , 
        \MSS_ADLIB_INST_GPOE[12] , \MSS_ADLIB_INST_GPOE[11] , 
        \MSS_ADLIB_INST_GPOE[10] , \MSS_ADLIB_INST_GPOE[9] , 
        \MSS_ADLIB_INST_GPOE[8] , \MSS_ADLIB_INST_GPOE[7] , 
        \MSS_ADLIB_INST_GPOE[6] , \MSS_ADLIB_INST_GPOE[5] , 
        \MSS_ADLIB_INST_GPOE[4] , \MSS_ADLIB_INST_GPOE[3] , 
        \MSS_ADLIB_INST_GPOE[2] , \MSS_ADLIB_INST_GPOE[1] , 
        \MSS_ADLIB_INST_GPOE[0] }), .SPI0DO(MSS_ADLIB_INST_SPI0DO), 
        .SPI0DOE(MSS_ADLIB_INST_SPI0DOE), .SPI0DI(crc_ahb_ip_MSS_GND), 
        .SPI0CLKI(crc_ahb_ip_MSS_GND), .SPI0CLKO(
        MSS_ADLIB_INST_SPI0CLKO), .SPI0MODE(MSS_ADLIB_INST_SPI0MODE), 
        .SPI0SSI(crc_ahb_ip_MSS_GND), .SPI0SSO({
        \MSS_ADLIB_INST_SPI0SSO[7] , \MSS_ADLIB_INST_SPI0SSO[6] , 
        \MSS_ADLIB_INST_SPI0SSO[5] , \MSS_ADLIB_INST_SPI0SSO[4] , 
        \MSS_ADLIB_INST_SPI0SSO[3] , \MSS_ADLIB_INST_SPI0SSO[2] , 
        \MSS_ADLIB_INST_SPI0SSO[1] , \MSS_ADLIB_INST_SPI0SSO[0] }), 
        .UART0TXD(MSS_UART_0_TXD_D), .UART0RXD(MSS_UART_0_RXD_Y), 
        .I2C0SDAI(crc_ahb_ip_MSS_GND), .I2C0SDAO(
        MSS_ADLIB_INST_I2C0SDAO), .I2C0SCLI(crc_ahb_ip_MSS_GND), 
        .I2C0SCLO(MSS_ADLIB_INST_I2C0SCLO), .SPI1DO(
        MSS_ADLIB_INST_SPI1DO), .SPI1DOE(MSS_ADLIB_INST_SPI1DOE), 
        .SPI1DI(crc_ahb_ip_MSS_GND), .SPI1CLKI(crc_ahb_ip_MSS_GND), 
        .SPI1CLKO(MSS_ADLIB_INST_SPI1CLKO), .SPI1MODE(
        MSS_ADLIB_INST_SPI1MODE), .SPI1SSI(crc_ahb_ip_MSS_GND), 
        .SPI1SSO({\MSS_ADLIB_INST_SPI1SSO[7] , 
        \MSS_ADLIB_INST_SPI1SSO[6] , \MSS_ADLIB_INST_SPI1SSO[5] , 
        \MSS_ADLIB_INST_SPI1SSO[4] , \MSS_ADLIB_INST_SPI1SSO[3] , 
        \MSS_ADLIB_INST_SPI1SSO[2] , \MSS_ADLIB_INST_SPI1SSO[1] , 
        \MSS_ADLIB_INST_SPI1SSO[0] }), .UART1TXD(
        MSS_ADLIB_INST_UART1TXD), .UART1RXD(crc_ahb_ip_MSS_GND), 
        .I2C1SDAI(crc_ahb_ip_MSS_GND), .I2C1SDAO(
        MSS_ADLIB_INST_I2C1SDAO), .I2C1SCLI(crc_ahb_ip_MSS_GND), 
        .I2C1SCLO(MSS_ADLIB_INST_I2C1SCLO), .MACTXD({
        \MSS_ADLIB_INST_MACTXD[1] , \MSS_ADLIB_INST_MACTXD[0] }), 
        .MACRXD({crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND}), .MACTXEN(
        MSS_ADLIB_INST_MACTXEN), .MACCRSDV(crc_ahb_ip_MSS_GND), 
        .MACRXER(crc_ahb_ip_MSS_GND), .MACMDI(crc_ahb_ip_MSS_GND), 
        .MACMDO(MSS_ADLIB_INST_MACMDO), .MACMDEN(
        MSS_ADLIB_INST_MACMDEN), .MACMDC(MSS_ADLIB_INST_MACMDC), 
        .EMCCLK(MSS_ADLIB_INST_EMCCLK), .EMCCLKRTN(
        MSS_ADLIB_INST_EMCCLK), .EMCRDB({crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, 
        crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND, crc_ahb_ip_MSS_GND}), 
        .EMCAB({\MSS_ADLIB_INST_EMCAB[25] , \MSS_ADLIB_INST_EMCAB[24] , 
        \MSS_ADLIB_INST_EMCAB[23] , \MSS_ADLIB_INST_EMCAB[22] , 
        \MSS_ADLIB_INST_EMCAB[21] , \MSS_ADLIB_INST_EMCAB[20] , 
        \MSS_ADLIB_INST_EMCAB[19] , \MSS_ADLIB_INST_EMCAB[18] , 
        \MSS_ADLIB_INST_EMCAB[17] , \MSS_ADLIB_INST_EMCAB[16] , 
        \MSS_ADLIB_INST_EMCAB[15] , \MSS_ADLIB_INST_EMCAB[14] , 
        \MSS_ADLIB_INST_EMCAB[13] , \MSS_ADLIB_INST_EMCAB[12] , 
        \MSS_ADLIB_INST_EMCAB[11] , \MSS_ADLIB_INST_EMCAB[10] , 
        \MSS_ADLIB_INST_EMCAB[9] , \MSS_ADLIB_INST_EMCAB[8] , 
        \MSS_ADLIB_INST_EMCAB[7] , \MSS_ADLIB_INST_EMCAB[6] , 
        \MSS_ADLIB_INST_EMCAB[5] , \MSS_ADLIB_INST_EMCAB[4] , 
        \MSS_ADLIB_INST_EMCAB[3] , \MSS_ADLIB_INST_EMCAB[2] , 
        \MSS_ADLIB_INST_EMCAB[1] , \MSS_ADLIB_INST_EMCAB[0] }), 
        .EMCWDB({\MSS_ADLIB_INST_EMCWDB[15] , 
        \MSS_ADLIB_INST_EMCWDB[14] , \MSS_ADLIB_INST_EMCWDB[13] , 
        \MSS_ADLIB_INST_EMCWDB[12] , \MSS_ADLIB_INST_EMCWDB[11] , 
        \MSS_ADLIB_INST_EMCWDB[10] , \MSS_ADLIB_INST_EMCWDB[9] , 
        \MSS_ADLIB_INST_EMCWDB[8] , \MSS_ADLIB_INST_EMCWDB[7] , 
        \MSS_ADLIB_INST_EMCWDB[6] , \MSS_ADLIB_INST_EMCWDB[5] , 
        \MSS_ADLIB_INST_EMCWDB[4] , \MSS_ADLIB_INST_EMCWDB[3] , 
        \MSS_ADLIB_INST_EMCWDB[2] , \MSS_ADLIB_INST_EMCWDB[1] , 
        \MSS_ADLIB_INST_EMCWDB[0] }), .EMCRWn(MSS_ADLIB_INST_EMCRWn), 
        .EMCCS0n(MSS_ADLIB_INST_EMCCS0n), .EMCCS1n(
        MSS_ADLIB_INST_EMCCS1n), .EMCOEN0n(MSS_ADLIB_INST_EMCOEN0n), 
        .EMCOEN1n(MSS_ADLIB_INST_EMCOEN1n), .EMCBYTEN({
        \MSS_ADLIB_INST_EMCBYTEN[1] , \MSS_ADLIB_INST_EMCBYTEN[0] }), 
        .EMCDBOE(MSS_ADLIB_INST_EMCDBOE), .ADC0(crc_ahb_ip_MSS_GND), 
        .ADC1(crc_ahb_ip_MSS_GND), .ADC2(crc_ahb_ip_MSS_GND), .ADC3(
        crc_ahb_ip_MSS_GND), .ADC4(crc_ahb_ip_MSS_GND), .ADC5(
        crc_ahb_ip_MSS_GND), .ADC6(crc_ahb_ip_MSS_GND), .ADC7(
        crc_ahb_ip_MSS_GND), .ADC8(crc_ahb_ip_MSS_GND), .ADC9(
        crc_ahb_ip_MSS_GND), .ADC10(crc_ahb_ip_MSS_GND), .ADC11(
        crc_ahb_ip_MSS_GND), .SDD0(MSS_ADLIB_INST_SDD0), .SDD1(
        MSS_ADLIB_INST_SDD1), .SDD2(MSS_ADLIB_INST_SDD2), .ABPS0(
        crc_ahb_ip_MSS_GND), .ABPS1(crc_ahb_ip_MSS_GND), .ABPS2(
        crc_ahb_ip_MSS_GND), .ABPS3(crc_ahb_ip_MSS_GND), .ABPS4(
        crc_ahb_ip_MSS_GND), .ABPS5(crc_ahb_ip_MSS_GND), .ABPS6(
        crc_ahb_ip_MSS_GND), .ABPS7(crc_ahb_ip_MSS_GND), .ABPS8(
        crc_ahb_ip_MSS_GND), .ABPS9(crc_ahb_ip_MSS_GND), .ABPS10(
        crc_ahb_ip_MSS_GND), .ABPS11(crc_ahb_ip_MSS_GND), .TM0(
        crc_ahb_ip_MSS_GND), .TM1(crc_ahb_ip_MSS_GND), .TM2(
        crc_ahb_ip_MSS_GND), .TM3(crc_ahb_ip_MSS_GND), .TM4(
        crc_ahb_ip_MSS_GND), .TM5(crc_ahb_ip_MSS_GND), .CM0(
        crc_ahb_ip_MSS_GND), .CM1(crc_ahb_ip_MSS_GND), .CM2(
        crc_ahb_ip_MSS_GND), .CM3(crc_ahb_ip_MSS_GND), .CM4(
        crc_ahb_ip_MSS_GND), .CM5(crc_ahb_ip_MSS_GND), .GNDTM0(
        crc_ahb_ip_MSS_GND), .GNDTM1(crc_ahb_ip_MSS_GND), .GNDTM2(
        crc_ahb_ip_MSS_GND), .VAREF0(crc_ahb_ip_MSS_GND), .VAREF1(
        crc_ahb_ip_MSS_GND), .VAREF2(crc_ahb_ip_MSS_GND), .VAREFOUT(
        MSS_ADLIB_INST_VAREFOUT), .GNDVAREF(crc_ahb_ip_MSS_GND), .PUn(
        crc_ahb_ip_MSS_GND));
    VCC VCC_i (.Y(crc_ahb_ip_MSS_VCC));
    INBUF_MSS #( .ACT_CONFIG(0), .ACT_PIN("U18") )  MSS_UART_0_RXD (
        .PAD(UART_0_RXD), .Y(MSS_UART_0_RXD_Y));
    GND GND_i (.Y(crc_ahb_ip_MSS_GND));
    
endmodule


module crc_ahb_ip(
       MSS_RESET_N,
       UART_0_RXD,
       UART_0_TXD
    );
input  MSS_RESET_N;
input  UART_0_RXD;
output UART_0_TXD;

    wire FAB_CLK, crc_ahb_ip_MSS_0_M2F_RESET_N, 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[2] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[3] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[4] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[16] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[17] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[18] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[19] , GND, 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK, 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[0] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS[1] , 
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE, 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[0] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[2] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[3] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[4] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[5] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[6] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[7] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[8] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[9] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[10] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[11] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[12] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[13] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[14] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[15] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[16] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[17] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[18] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[19] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[20] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[21] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[22] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[23] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[24] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[25] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[26] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[27] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[28] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[29] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[30] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[31] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[0] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[2] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[3] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[4] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[5] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[6] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[7] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[8] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[9] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[10] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[11] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[12] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[13] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[14] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[15] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[16] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[17] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[18] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[19] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[20] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[21] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[22] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[23] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[24] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[25] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[26] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[27] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[28] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[29] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[30] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[31] , VCC, N_153, 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[20] , N_363, N_355, 
        \crc_ip_0.CRC_UNIT.DATAPATH.crc_poly_size_77 , N_354, 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[19] , N_333, N_362, 
        \crc_ip_0.bus_wr[3] , N_365, \crc_ip_0.bus_wr[25] , N_336, 
        N_360, N_352, \crc_ip_0.bus_wr[1] , N_357, N_332, N_340, N_341, 
        N_342, N_387, N_5, CoreAHBLite_0_AHBmslave5_HREADY_i_0, N_347, 
        \crc_ip_0.bus_wr[0] , N_350, 
        \CoreAHBLite_0.matrix4x16.slavestage_5.un1_masterAddrInProg_6 , 
        \crc_ip_0.bus_wr[2] , N_349, N_348, 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[25] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[8] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[24] , N_351, N_367, 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[11] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[12] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[13] , N_356, N_361, 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[14] , N_358, N_366, 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[9] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[10] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[15] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[16] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[17] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[18] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[21] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[22] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[23] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[26] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[27] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[28] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[29] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[30] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[31] , N_364, 
        \crc_ip_0.bus_wr[16] , N_353, N_337, N_335, N_334, N_409, 
        N_408, \crc_ip_0.HOST_INTERFACE.HRDATA_0[23] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[22] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[21] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[18] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[1] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[1] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[5] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[5] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[3] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[3] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[10] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[9] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[8] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[24] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[25] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[27] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[7] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[7] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[13] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[4] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[4] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[19] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[14] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[30] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[16] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[12] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[11] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[26] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[29] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[28] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[0] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[0] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[6] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[6] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[17] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[2] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[2] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[31] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[15] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[20] , 
        defSlaveSMCurrentState_RNI5UNRI, crc_poly_size_77;
    
    CLKINT I_131 (.A(crc_poly_size_77), .Y(
        \crc_ip_0.CRC_UNIT.DATAPATH.crc_poly_size_77 ));
    CoreAHBLite_Z3 CoreAHBLite_0 (
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS({
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS[1] }), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE({
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[0] }), .HRDATA_2({
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[7] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[6] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[5] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[4] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[3] }), .HRDATA_1({
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[7] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[6] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[5] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[4] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[3] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[2] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[1] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[0] }), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_15(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[17] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_14(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[16] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[18] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[19] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[4] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_1(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[3] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_0(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[2] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA({
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[31] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[30] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[29] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[28] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[27] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[26] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[25] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[24] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[23] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[22] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[21] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[20] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[19] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[18] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[17] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[16] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[15] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[14] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[13] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[12] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[11] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[10] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[9] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[8] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[7] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[6] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[5] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[4] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[3] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[2] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[0] }), 
        .un4_HRDATA({\crc_ip_0.HOST_INTERFACE.un4_HRDATA[31] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[30] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[29] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[28] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[27] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[26] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[25] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[24] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[23] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[22] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[21] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[20] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[19] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[18] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[17] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[16] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[15] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[14] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[13] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[12] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[11] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[10] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[9] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[8] }), .HRDATA_0_1(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[1] ), .HRDATA_0_9(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[9] ), .HRDATA_0_10(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[10] ), .HRDATA_0_15(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[15] ), .HRDATA_0_16(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[16] ), .HRDATA_0_17(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[17] ), .HRDATA_0_18(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[18] ), .HRDATA_0_21(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[21] ), .HRDATA_0_22(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[22] ), .HRDATA_0_23(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[23] ), .HRDATA_0_26(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[26] ), .HRDATA_0_27(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[27] ), .HRDATA_0_28(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[28] ), .HRDATA_0_29(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[29] ), .HRDATA_0_30(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[30] ), .HRDATA_0_31(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[31] ), .HRDATA_0_14(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[14] ), .HRDATA_0_13(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[13] ), .HRDATA_0_12(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[12] ), .HRDATA_0_11(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[11] ), .HRDATA_0_24(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[24] ), .HRDATA_0_8(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[8] ), .HRDATA_0_25(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[25] ), .HRDATA_0_2(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[2] ), .HRDATA_0_0(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[0] ), .HRDATA_0_19(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[19] ), .HRDATA_0_20(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[20] ), .bus_wr_25(
        \crc_ip_0.bus_wr[25] ), .bus_wr_0(\crc_ip_0.bus_wr[0] ), 
        .bus_wr_1(\crc_ip_0.bus_wr[1] ), .bus_wr_2(
        \crc_ip_0.bus_wr[2] ), .bus_wr_16(\crc_ip_0.bus_wr[16] ), 
        .bus_wr_3(\crc_ip_0.bus_wr[3] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA({
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[31] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[30] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[29] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[28] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[27] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[26] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[25] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[24] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[23] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[22] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[21] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[20] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[19] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[18] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[17] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[16] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[15] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[14] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[13] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[12] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[11] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[10] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[9] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[8] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[7] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[6] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[5] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[4] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[3] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[2] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[0] }), 
        .defSlaveSMCurrentState_RNI5UNRI(
        defSlaveSMCurrentState_RNI5UNRI), 
        .CoreAHBLite_0_AHBmslave5_HREADY_i_0(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK), .N_153(N_153), 
        .FAB_CLK(FAB_CLK), .crc_ahb_ip_MSS_0_M2F_RESET_N(
        crc_ahb_ip_MSS_0_M2F_RESET_N), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE), .N_332(N_332), 
        .N_333(N_333), .N_334(N_334), .N_335(N_335), .N_336(N_336), 
        .N_337(N_337), .N_347(N_347), .N_348(N_348), .N_352(N_352), 
        .N_353(N_353), .N_358(N_358), .N_360(N_360), .N_361(N_361), 
        .N_364(N_364), .N_365(N_365), .N_366(N_366), .N_367(N_367), 
        .N_350(N_350), .N_357(N_357), .N_356(N_356), .N_351(N_351), 
        .N_349(N_349), .N_354(N_354), .N_362(N_362), .N_355(N_355), 
        .N_363(N_363), .un1_masterAddrInProg_6(
        \CoreAHBLite_0.matrix4x16.slavestage_5.un1_masterAddrInProg_6 )
        , .N_387(N_387), .N_408(N_408), .N_409(N_409), .N_5(N_5), 
        .N_342(N_342), .N_341(N_341), .N_340(N_340));
    crc_ip crc_ip_0 (.HRDATA_2({\crc_ip_0.HOST_INTERFACE.HRDATA_2[7] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[6] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[5] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[4] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_2[3] }), .HRDATA_1({
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[7] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[6] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[5] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[4] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[3] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[2] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[1] , 
        \crc_ip_0.HOST_INTERFACE.HRDATA_1[0] }), .HRDATA_0_20(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[20] ), .HRDATA_0_15(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[15] ), .HRDATA_0_31(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[31] ), .HRDATA_0_2(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[2] ), .HRDATA_0_17(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[17] ), .HRDATA_0_0(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[0] ), .HRDATA_0_28(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[28] ), .HRDATA_0_29(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[29] ), .HRDATA_0_26(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[26] ), .HRDATA_0_11(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[11] ), .HRDATA_0_12(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[12] ), .HRDATA_0_16(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[16] ), .HRDATA_0_30(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[30] ), .HRDATA_0_14(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[14] ), .HRDATA_0_19(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[19] ), .HRDATA_0_13(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[13] ), .HRDATA_0_27(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[27] ), .HRDATA_0_25(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[25] ), .HRDATA_0_24(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[24] ), .HRDATA_0_8(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[8] ), .HRDATA_0_9(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[9] ), .HRDATA_0_10(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[10] ), .HRDATA_0_1(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[1] ), .HRDATA_0_18(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[18] ), .HRDATA_0_21(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[21] ), .HRDATA_0_22(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[22] ), .HRDATA_0_23(
        \crc_ip_0.HOST_INTERFACE.HRDATA_0[23] ), .un4_HRDATA({
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[31] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[30] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[29] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[28] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[27] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[26] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[25] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[24] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[23] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[22] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[21] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[20] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[19] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[18] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[17] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[16] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[15] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[14] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[13] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[12] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[11] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[10] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[9] , 
        \crc_ip_0.HOST_INTERFACE.un4_HRDATA[8] }), .bus_wr_0(
        \crc_ip_0.bus_wr[0] ), .bus_wr_3(\crc_ip_0.bus_wr[3] ), 
        .bus_wr_1(\crc_ip_0.bus_wr[1] ), .bus_wr_16(
        \crc_ip_0.bus_wr[16] ), .bus_wr_25(\crc_ip_0.bus_wr[25] ), 
        .bus_wr_2(\crc_ip_0.bus_wr[2] ), .FAB_CLK(FAB_CLK), 
        .CoreAHBLite_0_AHBmslave5_HREADY_i_0(
        CoreAHBLite_0_AHBmslave5_HREADY_i_0), .N_347(N_347), 
        .crc_ahb_ip_MSS_0_M2F_RESET_N(crc_ahb_ip_MSS_0_M2F_RESET_N), 
        .N_350(N_350), .N_348(N_348), .N_349(N_349), 
        .un1_masterAddrInProg_6(
        \CoreAHBLite_0.matrix4x16.slavestage_5.un1_masterAddrInProg_6 )
        , .N_5(N_5), .N_408(N_408), .N_409(N_409), .N_387(N_387), 
        .N_340(N_340), .N_341(N_341), .N_342(N_342), .N_352(N_352), 
        .N_353(N_353), .N_358(N_358), .N_360(N_360), .N_361(N_361), 
        .N_364(N_364), .N_365(N_365), .N_366(N_366), .N_332(N_332), 
        .N_333(N_333), .N_334(N_334), .N_335(N_335), .N_336(N_336), 
        .N_337(N_337), .N_367(N_367), .crc_poly_size_77(
        crc_poly_size_77), .N_357(N_357), .N_356(N_356), .N_354(N_354), 
        .N_351(N_351), .N_362(N_362), .N_355(N_355), .N_363(N_363), 
        .crc_poly_size_77_0(
        \crc_ip_0.CRC_UNIT.DATAPATH.crc_poly_size_77 ));
    crc_ahb_ip_MSS crc_ahb_ip_MSS_0 (
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS({
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HTRANS[1] }), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_2(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[2] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_3(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[3] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_4(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[4] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_16(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[16] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_17(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[17] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_18(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[18] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR_19(
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HADDR[19] ), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA({
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[31] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[30] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[29] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[28] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[27] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[26] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[25] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[24] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[23] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[22] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[21] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[20] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[19] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[18] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[17] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[16] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[15] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[14] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[13] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[12] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[11] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[10] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[9] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[8] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[7] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[6] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[5] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[4] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[3] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[2] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWDATA[0] }), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA({
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[31] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[30] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[29] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[28] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[27] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[26] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[25] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[24] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[23] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[22] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[21] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[20] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[19] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[18] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[17] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[16] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[15] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[14] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[13] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[12] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[11] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[10] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[9] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[8] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[7] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[6] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[5] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[4] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[3] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[2] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HRDATA[0] }), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE({
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[1] , 
        \crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HSIZE[0] }), 
        .crc_ahb_ip_MSS_0_M2F_RESET_N(crc_ahb_ip_MSS_0_M2F_RESET_N), 
        .defSlaveSMCurrentState_RNI5UNRI(
        defSlaveSMCurrentState_RNI5UNRI), .UART_0_TXD(UART_0_TXD), 
        .UART_0_RXD(UART_0_RXD), .MSS_RESET_N(MSS_RESET_N), .FAB_CLK(
        FAB_CLK), .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HLOCK), 
        .crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE(
        crc_ahb_ip_MSS_0_MSS_MASTER_AHB_LITE_HWRITE), .N_153(N_153));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    
endmodule
